
module mem #(                   // 
    parameter  ADDR_LEN  = 11   // 
) (
    input  clk, rst,
    input  [ADDR_LEN-1:0] addr, // memory address
    output reg [31:0] rd_data,  // data read out
    input  wr_req,
    input  [31:0] wr_data       // data write in
);
localparam MEM_SIZE = 1<<ADDR_LEN;
reg [31:0] ram_cell [MEM_SIZE];

always @ (posedge clk or posedge rst)
    if(rst)
        rd_data <= 0;
    else
        rd_data <= ram_cell[addr];

always @ (posedge clk)
    if(wr_req) 
        ram_cell[addr] <= wr_data;

initial begin
    // dst matrix C
    ram_cell[       0] = 32'h0;  // 32'h225c5526;
    ram_cell[       1] = 32'h0;  // 32'hf4b4826b;
    ram_cell[       2] = 32'h0;  // 32'hbef276b4;
    ram_cell[       3] = 32'h0;  // 32'h290790ae;
    ram_cell[       4] = 32'h0;  // 32'h8c8db740;
    ram_cell[       5] = 32'h0;  // 32'h17248171;
    ram_cell[       6] = 32'h0;  // 32'had78d8f7;
    ram_cell[       7] = 32'h0;  // 32'h7b446b22;
    ram_cell[       8] = 32'h0;  // 32'hc04f049f;
    ram_cell[       9] = 32'h0;  // 32'hb7b52efc;
    ram_cell[      10] = 32'h0;  // 32'hd60fc807;
    ram_cell[      11] = 32'h0;  // 32'h303a1c37;
    ram_cell[      12] = 32'h0;  // 32'h1931cd11;
    ram_cell[      13] = 32'h0;  // 32'h171bc045;
    ram_cell[      14] = 32'h0;  // 32'h8892c914;
    ram_cell[      15] = 32'h0;  // 32'hd775026c;
    ram_cell[      16] = 32'h0;  // 32'ha02d0ca4;
    ram_cell[      17] = 32'h0;  // 32'hb4079d82;
    ram_cell[      18] = 32'h0;  // 32'he0b535d6;
    ram_cell[      19] = 32'h0;  // 32'h391bf2ca;
    ram_cell[      20] = 32'h0;  // 32'h90011639;
    ram_cell[      21] = 32'h0;  // 32'h496fa43c;
    ram_cell[      22] = 32'h0;  // 32'h83fea6a7;
    ram_cell[      23] = 32'h0;  // 32'hbd29893b;
    ram_cell[      24] = 32'h0;  // 32'h856ee5eb;
    ram_cell[      25] = 32'h0;  // 32'h91a256bf;
    ram_cell[      26] = 32'h0;  // 32'h673464ee;
    ram_cell[      27] = 32'h0;  // 32'h4aca6eb0;
    ram_cell[      28] = 32'h0;  // 32'ha5db0846;
    ram_cell[      29] = 32'h0;  // 32'h1c9838d2;
    ram_cell[      30] = 32'h0;  // 32'hde5adc2a;
    ram_cell[      31] = 32'h0;  // 32'h2eef9379;
    ram_cell[      32] = 32'h0;  // 32'h004b5ec4;
    ram_cell[      33] = 32'h0;  // 32'hc01ed742;
    ram_cell[      34] = 32'h0;  // 32'hc7b0719a;
    ram_cell[      35] = 32'h0;  // 32'h197eb23d;
    ram_cell[      36] = 32'h0;  // 32'hde198aa0;
    ram_cell[      37] = 32'h0;  // 32'h5cf7766e;
    ram_cell[      38] = 32'h0;  // 32'he3491734;
    ram_cell[      39] = 32'h0;  // 32'h3eb6b741;
    ram_cell[      40] = 32'h0;  // 32'he4a2197a;
    ram_cell[      41] = 32'h0;  // 32'h7e3d087d;
    ram_cell[      42] = 32'h0;  // 32'h7b9d9c2d;
    ram_cell[      43] = 32'h0;  // 32'h1f59bc99;
    ram_cell[      44] = 32'h0;  // 32'hd581e8ac;
    ram_cell[      45] = 32'h0;  // 32'hebf745a6;
    ram_cell[      46] = 32'h0;  // 32'h698e4fba;
    ram_cell[      47] = 32'h0;  // 32'h80f3d002;
    ram_cell[      48] = 32'h0;  // 32'h9eb3740f;
    ram_cell[      49] = 32'h0;  // 32'h8e67ba24;
    ram_cell[      50] = 32'h0;  // 32'h765ee8b7;
    ram_cell[      51] = 32'h0;  // 32'h0d93108d;
    ram_cell[      52] = 32'h0;  // 32'ha6a889a1;
    ram_cell[      53] = 32'h0;  // 32'h4dabfa66;
    ram_cell[      54] = 32'h0;  // 32'hc71c06d1;
    ram_cell[      55] = 32'h0;  // 32'h16f37e98;
    ram_cell[      56] = 32'h0;  // 32'h1fb75326;
    ram_cell[      57] = 32'h0;  // 32'he91725a2;
    ram_cell[      58] = 32'h0;  // 32'hadb6f493;
    ram_cell[      59] = 32'h0;  // 32'h6b7e8cff;
    ram_cell[      60] = 32'h0;  // 32'h27016aad;
    ram_cell[      61] = 32'h0;  // 32'hda059a4e;
    ram_cell[      62] = 32'h0;  // 32'h60fae404;
    ram_cell[      63] = 32'h0;  // 32'h2ae846f7;
    ram_cell[      64] = 32'h0;  // 32'h92017529;
    ram_cell[      65] = 32'h0;  // 32'h3aa37d85;
    ram_cell[      66] = 32'h0;  // 32'hd365ae88;
    ram_cell[      67] = 32'h0;  // 32'h77d6d49d;
    ram_cell[      68] = 32'h0;  // 32'h71e7f728;
    ram_cell[      69] = 32'h0;  // 32'h90a99089;
    ram_cell[      70] = 32'h0;  // 32'h1a3d3fb6;
    ram_cell[      71] = 32'h0;  // 32'h9eca312f;
    ram_cell[      72] = 32'h0;  // 32'h7e89a86b;
    ram_cell[      73] = 32'h0;  // 32'h859c8070;
    ram_cell[      74] = 32'h0;  // 32'h4b5d14ac;
    ram_cell[      75] = 32'h0;  // 32'h611e2af4;
    ram_cell[      76] = 32'h0;  // 32'h38be4f1f;
    ram_cell[      77] = 32'h0;  // 32'hed65e8b3;
    ram_cell[      78] = 32'h0;  // 32'h7b7ad5b5;
    ram_cell[      79] = 32'h0;  // 32'hba9f52fd;
    ram_cell[      80] = 32'h0;  // 32'h5f8e6a81;
    ram_cell[      81] = 32'h0;  // 32'h916bab8f;
    ram_cell[      82] = 32'h0;  // 32'heeaddace;
    ram_cell[      83] = 32'h0;  // 32'h739a97b8;
    ram_cell[      84] = 32'h0;  // 32'h9917facd;
    ram_cell[      85] = 32'h0;  // 32'hada8a1cc;
    ram_cell[      86] = 32'h0;  // 32'h7e6a1e34;
    ram_cell[      87] = 32'h0;  // 32'he18ce634;
    ram_cell[      88] = 32'h0;  // 32'he85f269c;
    ram_cell[      89] = 32'h0;  // 32'h7d903a02;
    ram_cell[      90] = 32'h0;  // 32'ha38afd80;
    ram_cell[      91] = 32'h0;  // 32'hfedb95d7;
    ram_cell[      92] = 32'h0;  // 32'hf8dc0888;
    ram_cell[      93] = 32'h0;  // 32'h05b0c206;
    ram_cell[      94] = 32'h0;  // 32'hc9921397;
    ram_cell[      95] = 32'h0;  // 32'hff238bd9;
    ram_cell[      96] = 32'h0;  // 32'hff783fab;
    ram_cell[      97] = 32'h0;  // 32'h87bee583;
    ram_cell[      98] = 32'h0;  // 32'h3b5696e1;
    ram_cell[      99] = 32'h0;  // 32'hec1852ae;
    ram_cell[     100] = 32'h0;  // 32'h1e6774ba;
    ram_cell[     101] = 32'h0;  // 32'h29ae4813;
    ram_cell[     102] = 32'h0;  // 32'he629bf2b;
    ram_cell[     103] = 32'h0;  // 32'h219254c1;
    ram_cell[     104] = 32'h0;  // 32'h34452942;
    ram_cell[     105] = 32'h0;  // 32'h0a36c48b;
    ram_cell[     106] = 32'h0;  // 32'h96318395;
    ram_cell[     107] = 32'h0;  // 32'h36e3f5e9;
    ram_cell[     108] = 32'h0;  // 32'hf28b36b9;
    ram_cell[     109] = 32'h0;  // 32'h3414299b;
    ram_cell[     110] = 32'h0;  // 32'h3d9082c4;
    ram_cell[     111] = 32'h0;  // 32'h99099d2d;
    ram_cell[     112] = 32'h0;  // 32'h7dd4f99d;
    ram_cell[     113] = 32'h0;  // 32'h50251729;
    ram_cell[     114] = 32'h0;  // 32'h6341e07a;
    ram_cell[     115] = 32'h0;  // 32'hafb0f975;
    ram_cell[     116] = 32'h0;  // 32'h5722cc9a;
    ram_cell[     117] = 32'h0;  // 32'hb61cd0b4;
    ram_cell[     118] = 32'h0;  // 32'hd34e3f9e;
    ram_cell[     119] = 32'h0;  // 32'h89f6a981;
    ram_cell[     120] = 32'h0;  // 32'he608f6bf;
    ram_cell[     121] = 32'h0;  // 32'he94eaf15;
    ram_cell[     122] = 32'h0;  // 32'hc52ea528;
    ram_cell[     123] = 32'h0;  // 32'h60c38c6e;
    ram_cell[     124] = 32'h0;  // 32'hc955709e;
    ram_cell[     125] = 32'h0;  // 32'h6592eda3;
    ram_cell[     126] = 32'h0;  // 32'h91bcfa28;
    ram_cell[     127] = 32'h0;  // 32'h73268867;
    ram_cell[     128] = 32'h0;  // 32'hfd811349;
    ram_cell[     129] = 32'h0;  // 32'hb4393eba;
    ram_cell[     130] = 32'h0;  // 32'h8b69cc10;
    ram_cell[     131] = 32'h0;  // 32'he62c300f;
    ram_cell[     132] = 32'h0;  // 32'h75f7dfcd;
    ram_cell[     133] = 32'h0;  // 32'h289bc546;
    ram_cell[     134] = 32'h0;  // 32'h83b5c155;
    ram_cell[     135] = 32'h0;  // 32'h1494f30d;
    ram_cell[     136] = 32'h0;  // 32'h0a16cebb;
    ram_cell[     137] = 32'h0;  // 32'h08f8a546;
    ram_cell[     138] = 32'h0;  // 32'hef348765;
    ram_cell[     139] = 32'h0;  // 32'h3833bc10;
    ram_cell[     140] = 32'h0;  // 32'hf370bab4;
    ram_cell[     141] = 32'h0;  // 32'h38ca7e1c;
    ram_cell[     142] = 32'h0;  // 32'hc2aa3cfc;
    ram_cell[     143] = 32'h0;  // 32'h4dbcbf05;
    ram_cell[     144] = 32'h0;  // 32'h4fc50c79;
    ram_cell[     145] = 32'h0;  // 32'h81c79f85;
    ram_cell[     146] = 32'h0;  // 32'haae8d9da;
    ram_cell[     147] = 32'h0;  // 32'ha6b93473;
    ram_cell[     148] = 32'h0;  // 32'h4cbc2e24;
    ram_cell[     149] = 32'h0;  // 32'haa1c1576;
    ram_cell[     150] = 32'h0;  // 32'hdf03e70a;
    ram_cell[     151] = 32'h0;  // 32'he1d6e0f9;
    ram_cell[     152] = 32'h0;  // 32'h421d6c0a;
    ram_cell[     153] = 32'h0;  // 32'hc02163b7;
    ram_cell[     154] = 32'h0;  // 32'h09716fa2;
    ram_cell[     155] = 32'h0;  // 32'h70adc72f;
    ram_cell[     156] = 32'h0;  // 32'hdd6a573e;
    ram_cell[     157] = 32'h0;  // 32'h8cdb7c3f;
    ram_cell[     158] = 32'h0;  // 32'hb18b8cf5;
    ram_cell[     159] = 32'h0;  // 32'h8804a79c;
    ram_cell[     160] = 32'h0;  // 32'ha412562d;
    ram_cell[     161] = 32'h0;  // 32'hd7379c17;
    ram_cell[     162] = 32'h0;  // 32'h37ffd5b9;
    ram_cell[     163] = 32'h0;  // 32'h95bb5cce;
    ram_cell[     164] = 32'h0;  // 32'h7b95a302;
    ram_cell[     165] = 32'h0;  // 32'h08342a60;
    ram_cell[     166] = 32'h0;  // 32'h5a50fedb;
    ram_cell[     167] = 32'h0;  // 32'h4e3719ff;
    ram_cell[     168] = 32'h0;  // 32'h66447920;
    ram_cell[     169] = 32'h0;  // 32'he24a4693;
    ram_cell[     170] = 32'h0;  // 32'h5d45c97d;
    ram_cell[     171] = 32'h0;  // 32'h240a864b;
    ram_cell[     172] = 32'h0;  // 32'h9ad20f38;
    ram_cell[     173] = 32'h0;  // 32'h45710b6d;
    ram_cell[     174] = 32'h0;  // 32'h26d380ef;
    ram_cell[     175] = 32'h0;  // 32'h776e6e89;
    ram_cell[     176] = 32'h0;  // 32'hc5e7d8ae;
    ram_cell[     177] = 32'h0;  // 32'h5e153a16;
    ram_cell[     178] = 32'h0;  // 32'h6d4e4466;
    ram_cell[     179] = 32'h0;  // 32'hac09d4fd;
    ram_cell[     180] = 32'h0;  // 32'hb6eb8c1d;
    ram_cell[     181] = 32'h0;  // 32'hb41fdb4f;
    ram_cell[     182] = 32'h0;  // 32'h32fbbf56;
    ram_cell[     183] = 32'h0;  // 32'h84e162b4;
    ram_cell[     184] = 32'h0;  // 32'h3d6a5302;
    ram_cell[     185] = 32'h0;  // 32'hb14d6a6a;
    ram_cell[     186] = 32'h0;  // 32'h2adb08df;
    ram_cell[     187] = 32'h0;  // 32'h1f896347;
    ram_cell[     188] = 32'h0;  // 32'hec00c32a;
    ram_cell[     189] = 32'h0;  // 32'h4b4c234d;
    ram_cell[     190] = 32'h0;  // 32'hd5103a4f;
    ram_cell[     191] = 32'h0;  // 32'h09749ca5;
    ram_cell[     192] = 32'h0;  // 32'h9b74fdb8;
    ram_cell[     193] = 32'h0;  // 32'h28d79bd1;
    ram_cell[     194] = 32'h0;  // 32'h46931389;
    ram_cell[     195] = 32'h0;  // 32'ha91d92a6;
    ram_cell[     196] = 32'h0;  // 32'hbc039e92;
    ram_cell[     197] = 32'h0;  // 32'habce0831;
    ram_cell[     198] = 32'h0;  // 32'h7cecf418;
    ram_cell[     199] = 32'h0;  // 32'hc2d7ca3a;
    ram_cell[     200] = 32'h0;  // 32'h1832897c;
    ram_cell[     201] = 32'h0;  // 32'hcfb79f53;
    ram_cell[     202] = 32'h0;  // 32'h99f24322;
    ram_cell[     203] = 32'h0;  // 32'h71c67295;
    ram_cell[     204] = 32'h0;  // 32'h518cf2e6;
    ram_cell[     205] = 32'h0;  // 32'hdc316970;
    ram_cell[     206] = 32'h0;  // 32'hb280f737;
    ram_cell[     207] = 32'h0;  // 32'h5877efc0;
    ram_cell[     208] = 32'h0;  // 32'hb6638b27;
    ram_cell[     209] = 32'h0;  // 32'h181c3814;
    ram_cell[     210] = 32'h0;  // 32'h14abc17a;
    ram_cell[     211] = 32'h0;  // 32'hb6cf66ba;
    ram_cell[     212] = 32'h0;  // 32'h7b9a955e;
    ram_cell[     213] = 32'h0;  // 32'hf9e87f99;
    ram_cell[     214] = 32'h0;  // 32'ha1b26783;
    ram_cell[     215] = 32'h0;  // 32'h2b2fb4ef;
    ram_cell[     216] = 32'h0;  // 32'h45e92693;
    ram_cell[     217] = 32'h0;  // 32'hac1f08a1;
    ram_cell[     218] = 32'h0;  // 32'hb9457ab5;
    ram_cell[     219] = 32'h0;  // 32'h54e70d82;
    ram_cell[     220] = 32'h0;  // 32'h2e99caff;
    ram_cell[     221] = 32'h0;  // 32'hc07bbc2e;
    ram_cell[     222] = 32'h0;  // 32'h2a3411ad;
    ram_cell[     223] = 32'h0;  // 32'hfffbcf12;
    ram_cell[     224] = 32'h0;  // 32'hf0f77a70;
    ram_cell[     225] = 32'h0;  // 32'h983ea5bc;
    ram_cell[     226] = 32'h0;  // 32'h28a799be;
    ram_cell[     227] = 32'h0;  // 32'h8304df72;
    ram_cell[     228] = 32'h0;  // 32'h88bcc55b;
    ram_cell[     229] = 32'h0;  // 32'h184f01b6;
    ram_cell[     230] = 32'h0;  // 32'had65463e;
    ram_cell[     231] = 32'h0;  // 32'h11f61c6a;
    ram_cell[     232] = 32'h0;  // 32'h3a0c0e02;
    ram_cell[     233] = 32'h0;  // 32'h713e1838;
    ram_cell[     234] = 32'h0;  // 32'h912b0a35;
    ram_cell[     235] = 32'h0;  // 32'h16b70d40;
    ram_cell[     236] = 32'h0;  // 32'h48a9b5d9;
    ram_cell[     237] = 32'h0;  // 32'h87b62753;
    ram_cell[     238] = 32'h0;  // 32'h693aa394;
    ram_cell[     239] = 32'h0;  // 32'hb211aa89;
    ram_cell[     240] = 32'h0;  // 32'h8a370acb;
    ram_cell[     241] = 32'h0;  // 32'ha56e1e8d;
    ram_cell[     242] = 32'h0;  // 32'h43ada732;
    ram_cell[     243] = 32'h0;  // 32'h47c5c65f;
    ram_cell[     244] = 32'h0;  // 32'h909160a4;
    ram_cell[     245] = 32'h0;  // 32'h0c7a7b10;
    ram_cell[     246] = 32'h0;  // 32'h9b29f18a;
    ram_cell[     247] = 32'h0;  // 32'h10ca6c59;
    ram_cell[     248] = 32'h0;  // 32'h8e580d73;
    ram_cell[     249] = 32'h0;  // 32'hbd860b41;
    ram_cell[     250] = 32'h0;  // 32'hce995f92;
    ram_cell[     251] = 32'h0;  // 32'h40b6d145;
    ram_cell[     252] = 32'h0;  // 32'h3db944c7;
    ram_cell[     253] = 32'h0;  // 32'h89ba536b;
    ram_cell[     254] = 32'h0;  // 32'h7b02c801;
    ram_cell[     255] = 32'h0;  // 32'hc616b7b2;
    // src matrix A
    ram_cell[     256] = 32'h7e55169f;
    ram_cell[     257] = 32'h12fc479a;
    ram_cell[     258] = 32'h512024ab;
    ram_cell[     259] = 32'h0e0860a7;
    ram_cell[     260] = 32'ha7644272;
    ram_cell[     261] = 32'h7c5710bf;
    ram_cell[     262] = 32'hb2e50a7f;
    ram_cell[     263] = 32'h154888b1;
    ram_cell[     264] = 32'hcd4fa6c5;
    ram_cell[     265] = 32'h216357c8;
    ram_cell[     266] = 32'hf861f372;
    ram_cell[     267] = 32'h9aac746d;
    ram_cell[     268] = 32'h04a72231;
    ram_cell[     269] = 32'hebd398c8;
    ram_cell[     270] = 32'h75c8b752;
    ram_cell[     271] = 32'h5c704ab8;
    ram_cell[     272] = 32'h45273a23;
    ram_cell[     273] = 32'hc2a1f47c;
    ram_cell[     274] = 32'h2b1c2604;
    ram_cell[     275] = 32'h96684292;
    ram_cell[     276] = 32'hf9fce4dd;
    ram_cell[     277] = 32'ha53e166e;
    ram_cell[     278] = 32'hb98e9847;
    ram_cell[     279] = 32'he4b7ec4b;
    ram_cell[     280] = 32'ha9c37ac7;
    ram_cell[     281] = 32'ha96ec8ba;
    ram_cell[     282] = 32'hab670245;
    ram_cell[     283] = 32'h3a3e7b65;
    ram_cell[     284] = 32'h98082e03;
    ram_cell[     285] = 32'h1cb2650d;
    ram_cell[     286] = 32'h6837da2f;
    ram_cell[     287] = 32'h881fab99;
    ram_cell[     288] = 32'h593bbb44;
    ram_cell[     289] = 32'hf11e4ed4;
    ram_cell[     290] = 32'h70f16038;
    ram_cell[     291] = 32'h9adacc4a;
    ram_cell[     292] = 32'hfd10a19a;
    ram_cell[     293] = 32'h9dad4ce4;
    ram_cell[     294] = 32'h14cc7564;
    ram_cell[     295] = 32'he7701014;
    ram_cell[     296] = 32'h58e0e828;
    ram_cell[     297] = 32'h69a46ebe;
    ram_cell[     298] = 32'h414c62af;
    ram_cell[     299] = 32'h129468f7;
    ram_cell[     300] = 32'hb2db875d;
    ram_cell[     301] = 32'h07e94b69;
    ram_cell[     302] = 32'h0fcba5cc;
    ram_cell[     303] = 32'heb609ecb;
    ram_cell[     304] = 32'h67bdbe65;
    ram_cell[     305] = 32'hf81689de;
    ram_cell[     306] = 32'hfe4f73cd;
    ram_cell[     307] = 32'ha134e1e6;
    ram_cell[     308] = 32'h125c7fc6;
    ram_cell[     309] = 32'h064b6a81;
    ram_cell[     310] = 32'ha37d580c;
    ram_cell[     311] = 32'h84292840;
    ram_cell[     312] = 32'hbb8fe381;
    ram_cell[     313] = 32'hef49042f;
    ram_cell[     314] = 32'hc0560440;
    ram_cell[     315] = 32'h0079ce80;
    ram_cell[     316] = 32'h29bbf883;
    ram_cell[     317] = 32'h3c8a3691;
    ram_cell[     318] = 32'h04481bed;
    ram_cell[     319] = 32'h65f68730;
    ram_cell[     320] = 32'h94e76169;
    ram_cell[     321] = 32'hd2f3de83;
    ram_cell[     322] = 32'hb0010fda;
    ram_cell[     323] = 32'h60bc59b4;
    ram_cell[     324] = 32'h142eb4f8;
    ram_cell[     325] = 32'hb51831d4;
    ram_cell[     326] = 32'h764c21fb;
    ram_cell[     327] = 32'h70aa58fa;
    ram_cell[     328] = 32'hf301d260;
    ram_cell[     329] = 32'h37a941e2;
    ram_cell[     330] = 32'hdeb17040;
    ram_cell[     331] = 32'h064b4437;
    ram_cell[     332] = 32'h94c462e4;
    ram_cell[     333] = 32'hfa0c9f3f;
    ram_cell[     334] = 32'h0834c4da;
    ram_cell[     335] = 32'hc55a3bdf;
    ram_cell[     336] = 32'hd15755c6;
    ram_cell[     337] = 32'hb26a5be0;
    ram_cell[     338] = 32'hc8d8851c;
    ram_cell[     339] = 32'h9a0bef1a;
    ram_cell[     340] = 32'h2e252c05;
    ram_cell[     341] = 32'h44092ad6;
    ram_cell[     342] = 32'h8a8f27db;
    ram_cell[     343] = 32'hacb55682;
    ram_cell[     344] = 32'h68f62a11;
    ram_cell[     345] = 32'h5cc1f302;
    ram_cell[     346] = 32'h6b1be21a;
    ram_cell[     347] = 32'h0e88ebd9;
    ram_cell[     348] = 32'hb38f9817;
    ram_cell[     349] = 32'h5f5821c5;
    ram_cell[     350] = 32'ha5d20387;
    ram_cell[     351] = 32'h8c59f00c;
    ram_cell[     352] = 32'hc2eb3bfb;
    ram_cell[     353] = 32'hd65bebc1;
    ram_cell[     354] = 32'h99d5ad0b;
    ram_cell[     355] = 32'h25608690;
    ram_cell[     356] = 32'hb1d4f597;
    ram_cell[     357] = 32'hfffe08aa;
    ram_cell[     358] = 32'haf79784a;
    ram_cell[     359] = 32'h7fbd8ff5;
    ram_cell[     360] = 32'h8bbfa3ad;
    ram_cell[     361] = 32'h0e58252e;
    ram_cell[     362] = 32'h497c465d;
    ram_cell[     363] = 32'hc30b419d;
    ram_cell[     364] = 32'ha9fcb6b9;
    ram_cell[     365] = 32'h707ab218;
    ram_cell[     366] = 32'h0c222c9f;
    ram_cell[     367] = 32'had55bc45;
    ram_cell[     368] = 32'h4711f9a5;
    ram_cell[     369] = 32'h285a207f;
    ram_cell[     370] = 32'h51103abc;
    ram_cell[     371] = 32'h896eb00c;
    ram_cell[     372] = 32'h773a6be4;
    ram_cell[     373] = 32'h8ecbaf1b;
    ram_cell[     374] = 32'h531fb7ee;
    ram_cell[     375] = 32'hd6048165;
    ram_cell[     376] = 32'h52ebe2c7;
    ram_cell[     377] = 32'h6d5fc8ad;
    ram_cell[     378] = 32'h7cc6d209;
    ram_cell[     379] = 32'h30f9ab42;
    ram_cell[     380] = 32'h3a80b95e;
    ram_cell[     381] = 32'h0537e949;
    ram_cell[     382] = 32'hef427578;
    ram_cell[     383] = 32'h42ffe82f;
    ram_cell[     384] = 32'he86854f4;
    ram_cell[     385] = 32'h6ebbc846;
    ram_cell[     386] = 32'h6a3b0060;
    ram_cell[     387] = 32'hd762650f;
    ram_cell[     388] = 32'h2de5ecbf;
    ram_cell[     389] = 32'hb6f7a823;
    ram_cell[     390] = 32'h2ddb79df;
    ram_cell[     391] = 32'hc93b05e4;
    ram_cell[     392] = 32'hb991bd26;
    ram_cell[     393] = 32'h35908796;
    ram_cell[     394] = 32'h1ddf819b;
    ram_cell[     395] = 32'hd447f402;
    ram_cell[     396] = 32'h50fda332;
    ram_cell[     397] = 32'h24396b3b;
    ram_cell[     398] = 32'hf3c0a2ef;
    ram_cell[     399] = 32'ha5efa6cd;
    ram_cell[     400] = 32'h634f57d5;
    ram_cell[     401] = 32'h9dd63d5c;
    ram_cell[     402] = 32'h0881244c;
    ram_cell[     403] = 32'hb99cfd0f;
    ram_cell[     404] = 32'h32814b3c;
    ram_cell[     405] = 32'h67a5cda8;
    ram_cell[     406] = 32'h8dde5e39;
    ram_cell[     407] = 32'ha7352340;
    ram_cell[     408] = 32'ha73d79a8;
    ram_cell[     409] = 32'h220f349d;
    ram_cell[     410] = 32'h718bd5d6;
    ram_cell[     411] = 32'hb044510a;
    ram_cell[     412] = 32'hda529014;
    ram_cell[     413] = 32'hdd6be97e;
    ram_cell[     414] = 32'h4ed975d1;
    ram_cell[     415] = 32'h3ecd6b38;
    ram_cell[     416] = 32'h50e80621;
    ram_cell[     417] = 32'h0377aac7;
    ram_cell[     418] = 32'hb22f6874;
    ram_cell[     419] = 32'h9385dd2d;
    ram_cell[     420] = 32'h453aea63;
    ram_cell[     421] = 32'h2ddf9505;
    ram_cell[     422] = 32'hbcee48e0;
    ram_cell[     423] = 32'h8551641c;
    ram_cell[     424] = 32'h90244358;
    ram_cell[     425] = 32'hb8d0e57c;
    ram_cell[     426] = 32'h51393fc9;
    ram_cell[     427] = 32'h6b988cb5;
    ram_cell[     428] = 32'h2db4ef23;
    ram_cell[     429] = 32'h93331a6d;
    ram_cell[     430] = 32'h39713439;
    ram_cell[     431] = 32'h62edb5de;
    ram_cell[     432] = 32'h7a320b58;
    ram_cell[     433] = 32'hb29132a4;
    ram_cell[     434] = 32'hb27d8a39;
    ram_cell[     435] = 32'h35492bac;
    ram_cell[     436] = 32'h66b15cd5;
    ram_cell[     437] = 32'h2e57ac4d;
    ram_cell[     438] = 32'h0fb55f8a;
    ram_cell[     439] = 32'h779bac90;
    ram_cell[     440] = 32'hadb04e7c;
    ram_cell[     441] = 32'h00de4f3a;
    ram_cell[     442] = 32'hd1322d37;
    ram_cell[     443] = 32'h375adda2;
    ram_cell[     444] = 32'h177beb3e;
    ram_cell[     445] = 32'h8fcfbec8;
    ram_cell[     446] = 32'h3445b74a;
    ram_cell[     447] = 32'h48918208;
    ram_cell[     448] = 32'hdd2f558b;
    ram_cell[     449] = 32'haff03801;
    ram_cell[     450] = 32'h9f4fe534;
    ram_cell[     451] = 32'h031ff76c;
    ram_cell[     452] = 32'hfcc7753c;
    ram_cell[     453] = 32'h96ee118a;
    ram_cell[     454] = 32'hb3bd7902;
    ram_cell[     455] = 32'h2a724a7a;
    ram_cell[     456] = 32'hccfc9d45;
    ram_cell[     457] = 32'h744144c8;
    ram_cell[     458] = 32'he2c61564;
    ram_cell[     459] = 32'h3ebd1e4e;
    ram_cell[     460] = 32'h79d8a972;
    ram_cell[     461] = 32'h354cea18;
    ram_cell[     462] = 32'h621a5cb9;
    ram_cell[     463] = 32'h366ec03a;
    ram_cell[     464] = 32'h84529344;
    ram_cell[     465] = 32'h0ee35704;
    ram_cell[     466] = 32'hd70805b0;
    ram_cell[     467] = 32'hbc6a01f8;
    ram_cell[     468] = 32'h51dcf034;
    ram_cell[     469] = 32'h9551bfe3;
    ram_cell[     470] = 32'h2f3b5a74;
    ram_cell[     471] = 32'h89de8ff0;
    ram_cell[     472] = 32'hdddc7dfc;
    ram_cell[     473] = 32'h08a0f1f9;
    ram_cell[     474] = 32'hcd78e9ef;
    ram_cell[     475] = 32'h69533dd2;
    ram_cell[     476] = 32'hb4445464;
    ram_cell[     477] = 32'hffd923f3;
    ram_cell[     478] = 32'ha2f5f420;
    ram_cell[     479] = 32'h782c0782;
    ram_cell[     480] = 32'h960c0731;
    ram_cell[     481] = 32'hd70d2768;
    ram_cell[     482] = 32'h629e8ac4;
    ram_cell[     483] = 32'h147d8082;
    ram_cell[     484] = 32'h76a2d1ee;
    ram_cell[     485] = 32'hb2cfef29;
    ram_cell[     486] = 32'h888af48e;
    ram_cell[     487] = 32'he979ce82;
    ram_cell[     488] = 32'h27db6188;
    ram_cell[     489] = 32'h2ab68996;
    ram_cell[     490] = 32'h558880cb;
    ram_cell[     491] = 32'h2786ebc7;
    ram_cell[     492] = 32'hd649076f;
    ram_cell[     493] = 32'had0f6336;
    ram_cell[     494] = 32'hfa81183e;
    ram_cell[     495] = 32'h32eec9cb;
    ram_cell[     496] = 32'h41d54fe3;
    ram_cell[     497] = 32'h28f79e6e;
    ram_cell[     498] = 32'h1c3f41a3;
    ram_cell[     499] = 32'h284fbd24;
    ram_cell[     500] = 32'hf94ac77c;
    ram_cell[     501] = 32'h3d71d361;
    ram_cell[     502] = 32'he59e634f;
    ram_cell[     503] = 32'h2d5e80f3;
    ram_cell[     504] = 32'hb73db23c;
    ram_cell[     505] = 32'h7f79953c;
    ram_cell[     506] = 32'h70b7238b;
    ram_cell[     507] = 32'h9a1020bd;
    ram_cell[     508] = 32'h74e52727;
    ram_cell[     509] = 32'hfd9b1855;
    ram_cell[     510] = 32'hbf73b950;
    ram_cell[     511] = 32'hf2e25be9;
    // src matrix B
    ram_cell[     512] = 32'h248a622e;
    ram_cell[     513] = 32'hdbba9a63;
    ram_cell[     514] = 32'h932eb330;
    ram_cell[     515] = 32'hb83a0974;
    ram_cell[     516] = 32'hb976be73;
    ram_cell[     517] = 32'h181f3b26;
    ram_cell[     518] = 32'h1d59eac9;
    ram_cell[     519] = 32'hd82582f5;
    ram_cell[     520] = 32'hf2e0bbcf;
    ram_cell[     521] = 32'h04ad78fe;
    ram_cell[     522] = 32'hfb669d7d;
    ram_cell[     523] = 32'h70fb5830;
    ram_cell[     524] = 32'had48a36e;
    ram_cell[     525] = 32'hedc90170;
    ram_cell[     526] = 32'hd45f207d;
    ram_cell[     527] = 32'ha8f8b8f6;
    ram_cell[     528] = 32'h4f1a7ae4;
    ram_cell[     529] = 32'hdb589e97;
    ram_cell[     530] = 32'h599d00c1;
    ram_cell[     531] = 32'hb935d3de;
    ram_cell[     532] = 32'h5021b9ab;
    ram_cell[     533] = 32'h31bda760;
    ram_cell[     534] = 32'h77f314ca;
    ram_cell[     535] = 32'hbf6dc966;
    ram_cell[     536] = 32'h2670c4a0;
    ram_cell[     537] = 32'hfda6b2b5;
    ram_cell[     538] = 32'h2a3fc53a;
    ram_cell[     539] = 32'hebf280be;
    ram_cell[     540] = 32'h4148eff7;
    ram_cell[     541] = 32'habf86782;
    ram_cell[     542] = 32'h5331f444;
    ram_cell[     543] = 32'h4bf0e98c;
    ram_cell[     544] = 32'h0ad646dc;
    ram_cell[     545] = 32'hec18f2fb;
    ram_cell[     546] = 32'ha38b1588;
    ram_cell[     547] = 32'hafe6e14c;
    ram_cell[     548] = 32'h23dbb03f;
    ram_cell[     549] = 32'h42a91e07;
    ram_cell[     550] = 32'h6a3cf7cf;
    ram_cell[     551] = 32'h723af3d1;
    ram_cell[     552] = 32'h363e2f0e;
    ram_cell[     553] = 32'h56fe1ffc;
    ram_cell[     554] = 32'h9ef8dc79;
    ram_cell[     555] = 32'h24cb4bec;
    ram_cell[     556] = 32'h8bb0ee7b;
    ram_cell[     557] = 32'he4a3fada;
    ram_cell[     558] = 32'h1350326c;
    ram_cell[     559] = 32'h337aff1c;
    ram_cell[     560] = 32'h274a64e0;
    ram_cell[     561] = 32'hc496a0bd;
    ram_cell[     562] = 32'hfac7a47f;
    ram_cell[     563] = 32'h7675193a;
    ram_cell[     564] = 32'hb7dc2ea7;
    ram_cell[     565] = 32'hd91260eb;
    ram_cell[     566] = 32'h2ea635ea;
    ram_cell[     567] = 32'hbd608e66;
    ram_cell[     568] = 32'h2e516580;
    ram_cell[     569] = 32'h3596cd8e;
    ram_cell[     570] = 32'h51fc8bb4;
    ram_cell[     571] = 32'hedb2b30f;
    ram_cell[     572] = 32'hbd38a319;
    ram_cell[     573] = 32'h5077374c;
    ram_cell[     574] = 32'h38848c28;
    ram_cell[     575] = 32'h6d078c10;
    ram_cell[     576] = 32'h87e92831;
    ram_cell[     577] = 32'h98caa405;
    ram_cell[     578] = 32'h24ef16f6;
    ram_cell[     579] = 32'h97f9eb83;
    ram_cell[     580] = 32'hafc03c52;
    ram_cell[     581] = 32'h08573c68;
    ram_cell[     582] = 32'h402ca8a5;
    ram_cell[     583] = 32'h0f13581e;
    ram_cell[     584] = 32'h478acabe;
    ram_cell[     585] = 32'hd1413eeb;
    ram_cell[     586] = 32'h65287118;
    ram_cell[     587] = 32'hbb4b82cf;
    ram_cell[     588] = 32'h7b471431;
    ram_cell[     589] = 32'h8d5dde3c;
    ram_cell[     590] = 32'hc1731a00;
    ram_cell[     591] = 32'h4866fb7a;
    ram_cell[     592] = 32'hb25c1622;
    ram_cell[     593] = 32'h32099728;
    ram_cell[     594] = 32'h5d9ac432;
    ram_cell[     595] = 32'ha18e037c;
    ram_cell[     596] = 32'h2120def2;
    ram_cell[     597] = 32'h2a05bad4;
    ram_cell[     598] = 32'h7aefe8b4;
    ram_cell[     599] = 32'hcd643d52;
    ram_cell[     600] = 32'he838844b;
    ram_cell[     601] = 32'h880c322f;
    ram_cell[     602] = 32'h7e3e120a;
    ram_cell[     603] = 32'h10c76c07;
    ram_cell[     604] = 32'h7b1c8756;
    ram_cell[     605] = 32'hb4607297;
    ram_cell[     606] = 32'hd92af3f5;
    ram_cell[     607] = 32'h25771773;
    ram_cell[     608] = 32'h2f852b1d;
    ram_cell[     609] = 32'h2ad9f192;
    ram_cell[     610] = 32'ha1d9f71a;
    ram_cell[     611] = 32'h4aa56f6b;
    ram_cell[     612] = 32'h07b0988d;
    ram_cell[     613] = 32'h834e4988;
    ram_cell[     614] = 32'hf9297598;
    ram_cell[     615] = 32'h42b54ad7;
    ram_cell[     616] = 32'h25d173bb;
    ram_cell[     617] = 32'h93742df7;
    ram_cell[     618] = 32'h14d1ed03;
    ram_cell[     619] = 32'h63e63e25;
    ram_cell[     620] = 32'hb5402944;
    ram_cell[     621] = 32'h6fbb3ba1;
    ram_cell[     622] = 32'h24487e02;
    ram_cell[     623] = 32'h028cd0b0;
    ram_cell[     624] = 32'hf45bd2f4;
    ram_cell[     625] = 32'h601cb70b;
    ram_cell[     626] = 32'h77f13070;
    ram_cell[     627] = 32'hc680c33f;
    ram_cell[     628] = 32'h519e0921;
    ram_cell[     629] = 32'hb63e243d;
    ram_cell[     630] = 32'h7b7637e8;
    ram_cell[     631] = 32'hd697057b;
    ram_cell[     632] = 32'h520564aa;
    ram_cell[     633] = 32'hfa1901bc;
    ram_cell[     634] = 32'h9d0c6c08;
    ram_cell[     635] = 32'h9b84a50a;
    ram_cell[     636] = 32'hafbbf3f2;
    ram_cell[     637] = 32'h989fae07;
    ram_cell[     638] = 32'hd916b711;
    ram_cell[     639] = 32'hbc63c209;
    ram_cell[     640] = 32'h17dcc022;
    ram_cell[     641] = 32'ha1cae383;
    ram_cell[     642] = 32'hae011853;
    ram_cell[     643] = 32'h8449d015;
    ram_cell[     644] = 32'h180e7485;
    ram_cell[     645] = 32'h202cb61b;
    ram_cell[     646] = 32'h830e6928;
    ram_cell[     647] = 32'hca7ef4b6;
    ram_cell[     648] = 32'h7bcb08f4;
    ram_cell[     649] = 32'h9e488356;
    ram_cell[     650] = 32'h294e4d2f;
    ram_cell[     651] = 32'h1fa290e0;
    ram_cell[     652] = 32'ha73dc922;
    ram_cell[     653] = 32'hd6b008e5;
    ram_cell[     654] = 32'h1ec32216;
    ram_cell[     655] = 32'hee1357ff;
    ram_cell[     656] = 32'ha43eeb38;
    ram_cell[     657] = 32'ha7341ab7;
    ram_cell[     658] = 32'h6568f108;
    ram_cell[     659] = 32'habcca537;
    ram_cell[     660] = 32'heae80b70;
    ram_cell[     661] = 32'h45b0fb39;
    ram_cell[     662] = 32'hac1422a0;
    ram_cell[     663] = 32'h3afeea14;
    ram_cell[     664] = 32'hf56d6db7;
    ram_cell[     665] = 32'hd413b90e;
    ram_cell[     666] = 32'h221e85c2;
    ram_cell[     667] = 32'h82c46d62;
    ram_cell[     668] = 32'hcc381c04;
    ram_cell[     669] = 32'h9f548187;
    ram_cell[     670] = 32'h78f6c462;
    ram_cell[     671] = 32'hcb5ae46d;
    ram_cell[     672] = 32'h6c0c7d5d;
    ram_cell[     673] = 32'h203d2d9a;
    ram_cell[     674] = 32'hcde231b2;
    ram_cell[     675] = 32'h753658e0;
    ram_cell[     676] = 32'h390deabe;
    ram_cell[     677] = 32'h7f1aa7c4;
    ram_cell[     678] = 32'hd7153a76;
    ram_cell[     679] = 32'hbede7497;
    ram_cell[     680] = 32'h6ab6a15d;
    ram_cell[     681] = 32'h9bb95736;
    ram_cell[     682] = 32'h781f117e;
    ram_cell[     683] = 32'h52603679;
    ram_cell[     684] = 32'h5f458144;
    ram_cell[     685] = 32'hd06a48d6;
    ram_cell[     686] = 32'h6ce491c6;
    ram_cell[     687] = 32'h718bf260;
    ram_cell[     688] = 32'h6dd32ae2;
    ram_cell[     689] = 32'h55a909b7;
    ram_cell[     690] = 32'h025a4a51;
    ram_cell[     691] = 32'h2c9a17d6;
    ram_cell[     692] = 32'h5ef6596f;
    ram_cell[     693] = 32'he4afdaec;
    ram_cell[     694] = 32'h23eca0c2;
    ram_cell[     695] = 32'h770a6671;
    ram_cell[     696] = 32'h9b422b68;
    ram_cell[     697] = 32'hd0f33839;
    ram_cell[     698] = 32'h9284408c;
    ram_cell[     699] = 32'h6d16ae1d;
    ram_cell[     700] = 32'h0c1739f3;
    ram_cell[     701] = 32'hb39b0aff;
    ram_cell[     702] = 32'h1d4f0dd1;
    ram_cell[     703] = 32'h28b1af1a;
    ram_cell[     704] = 32'h4ba06d4b;
    ram_cell[     705] = 32'hac2266a7;
    ram_cell[     706] = 32'h14a635a1;
    ram_cell[     707] = 32'h0499f721;
    ram_cell[     708] = 32'h296258a3;
    ram_cell[     709] = 32'hf94bef1d;
    ram_cell[     710] = 32'h308f4afd;
    ram_cell[     711] = 32'hd975c49b;
    ram_cell[     712] = 32'h734eb146;
    ram_cell[     713] = 32'ha50476d7;
    ram_cell[     714] = 32'h254a774b;
    ram_cell[     715] = 32'hbf2a3711;
    ram_cell[     716] = 32'hf06c9948;
    ram_cell[     717] = 32'h146a4dda;
    ram_cell[     718] = 32'h900ec348;
    ram_cell[     719] = 32'h72a23791;
    ram_cell[     720] = 32'h1902ec9e;
    ram_cell[     721] = 32'h191b01cb;
    ram_cell[     722] = 32'h59cea6cc;
    ram_cell[     723] = 32'h5ecb9e15;
    ram_cell[     724] = 32'h7dfab2be;
    ram_cell[     725] = 32'h7da0942a;
    ram_cell[     726] = 32'h5625463b;
    ram_cell[     727] = 32'h5e063b6a;
    ram_cell[     728] = 32'hb81dd3f6;
    ram_cell[     729] = 32'he0a995c6;
    ram_cell[     730] = 32'hee4c6963;
    ram_cell[     731] = 32'hbf6b86da;
    ram_cell[     732] = 32'h64f0c65b;
    ram_cell[     733] = 32'hfac9e480;
    ram_cell[     734] = 32'h33daa542;
    ram_cell[     735] = 32'hc836b4f0;
    ram_cell[     736] = 32'h102a51a4;
    ram_cell[     737] = 32'h3e8e9f92;
    ram_cell[     738] = 32'h405edcd3;
    ram_cell[     739] = 32'he1c6bc2b;
    ram_cell[     740] = 32'h79061093;
    ram_cell[     741] = 32'hc8260b6a;
    ram_cell[     742] = 32'hb02f1139;
    ram_cell[     743] = 32'hb98fd875;
    ram_cell[     744] = 32'hb69b63bf;
    ram_cell[     745] = 32'hcb68f970;
    ram_cell[     746] = 32'h62408a42;
    ram_cell[     747] = 32'h6496dd23;
    ram_cell[     748] = 32'h0639b013;
    ram_cell[     749] = 32'h6a6d8d91;
    ram_cell[     750] = 32'h9f72476c;
    ram_cell[     751] = 32'h348ea3bb;
    ram_cell[     752] = 32'h59a83650;
    ram_cell[     753] = 32'hded2a95d;
    ram_cell[     754] = 32'h55e753d2;
    ram_cell[     755] = 32'hdf69bd33;
    ram_cell[     756] = 32'h0e2466c6;
    ram_cell[     757] = 32'h47c2cdcf;
    ram_cell[     758] = 32'h900083b4;
    ram_cell[     759] = 32'hbd2ff9d8;
    ram_cell[     760] = 32'he5483c65;
    ram_cell[     761] = 32'hcae86127;
    ram_cell[     762] = 32'h221c1267;
    ram_cell[     763] = 32'hf0081e5c;
    ram_cell[     764] = 32'h64ffc114;
    ram_cell[     765] = 32'h25498adb;
    ram_cell[     766] = 32'h1bc0c2e1;
    ram_cell[     767] = 32'h13f11619;
end

endmodule

