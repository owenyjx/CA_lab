    Usage:
        python generate_mem_for_quicksort.py [matrix size]
    Example:
        python generate_mem_for_quicksort.py 16
    Tip: use this command to write to file:
        python generate_mem_for_quicksort.py 16 > mem.sv
