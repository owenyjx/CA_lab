
module mem #(                   // 
    parameter  ADDR_LEN  = 11   // 
) (
    input  clk, rst,
    input  [ADDR_LEN-1:0] addr, // memory address
    output reg [31:0] rd_data,  // data read out
    input  wr_req,
    input  [31:0] wr_data       // data write in
);
localparam MEM_SIZE = 1<<ADDR_LEN;
reg [31:0] ram_cell [MEM_SIZE];

always @ (posedge clk or posedge rst)
    if(rst)
        rd_data <= 0;
    else
        rd_data <= ram_cell[addr];

always @ (posedge clk)
    if(wr_req) 
        ram_cell[addr] <= wr_data;

initial begin
    // dst matrix C
    ram_cell[       0] = 32'h0;  // 32'he956c8d3;
    ram_cell[       1] = 32'h0;  // 32'h06d96607;
    ram_cell[       2] = 32'h0;  // 32'hacca2120;
    ram_cell[       3] = 32'h0;  // 32'h32f8f3bb;
    ram_cell[       4] = 32'h0;  // 32'h74ff35a4;
    ram_cell[       5] = 32'h0;  // 32'hb1917463;
    ram_cell[       6] = 32'h0;  // 32'he4e069a7;
    ram_cell[       7] = 32'h0;  // 32'hd31685cb;
    ram_cell[       8] = 32'h0;  // 32'hf0292d2c;
    ram_cell[       9] = 32'h0;  // 32'h40ba8a1a;
    ram_cell[      10] = 32'h0;  // 32'h29b74833;
    ram_cell[      11] = 32'h0;  // 32'hfecbbb52;
    ram_cell[      12] = 32'h0;  // 32'ha9072aa4;
    ram_cell[      13] = 32'h0;  // 32'h40ab291a;
    ram_cell[      14] = 32'h0;  // 32'hc6edb65d;
    ram_cell[      15] = 32'h0;  // 32'h1f3225f1;
    ram_cell[      16] = 32'h0;  // 32'ha2fe9206;
    ram_cell[      17] = 32'h0;  // 32'h775a96d5;
    ram_cell[      18] = 32'h0;  // 32'hc58df6f5;
    ram_cell[      19] = 32'h0;  // 32'he234604e;
    ram_cell[      20] = 32'h0;  // 32'hafabc18d;
    ram_cell[      21] = 32'h0;  // 32'h4ba40c33;
    ram_cell[      22] = 32'h0;  // 32'hba5c9c6c;
    ram_cell[      23] = 32'h0;  // 32'h5992a322;
    ram_cell[      24] = 32'h0;  // 32'h03123710;
    ram_cell[      25] = 32'h0;  // 32'h058023c0;
    ram_cell[      26] = 32'h0;  // 32'h92237999;
    ram_cell[      27] = 32'h0;  // 32'ha7a0f62d;
    ram_cell[      28] = 32'h0;  // 32'h1d4819b2;
    ram_cell[      29] = 32'h0;  // 32'h5f64ca77;
    ram_cell[      30] = 32'h0;  // 32'h9efee40b;
    ram_cell[      31] = 32'h0;  // 32'h5e7c3910;
    ram_cell[      32] = 32'h0;  // 32'h70f1990b;
    ram_cell[      33] = 32'h0;  // 32'he76e3368;
    ram_cell[      34] = 32'h0;  // 32'hfa5e5027;
    ram_cell[      35] = 32'h0;  // 32'h955f9c61;
    ram_cell[      36] = 32'h0;  // 32'hfd5a285a;
    ram_cell[      37] = 32'h0;  // 32'h5d392731;
    ram_cell[      38] = 32'h0;  // 32'hc86da623;
    ram_cell[      39] = 32'h0;  // 32'hd181d540;
    ram_cell[      40] = 32'h0;  // 32'heae42e96;
    ram_cell[      41] = 32'h0;  // 32'hbd9dbbd3;
    ram_cell[      42] = 32'h0;  // 32'h348d1e24;
    ram_cell[      43] = 32'h0;  // 32'h53ced800;
    ram_cell[      44] = 32'h0;  // 32'hcf855fe8;
    ram_cell[      45] = 32'h0;  // 32'hbb53b919;
    ram_cell[      46] = 32'h0;  // 32'h0eae8fa5;
    ram_cell[      47] = 32'h0;  // 32'h048db3dc;
    ram_cell[      48] = 32'h0;  // 32'h9ad88810;
    ram_cell[      49] = 32'h0;  // 32'hfa3d0426;
    ram_cell[      50] = 32'h0;  // 32'h4993f6ce;
    ram_cell[      51] = 32'h0;  // 32'h3e6c7ad0;
    ram_cell[      52] = 32'h0;  // 32'h11ee4b63;
    ram_cell[      53] = 32'h0;  // 32'h4fd5b054;
    ram_cell[      54] = 32'h0;  // 32'hbac2859c;
    ram_cell[      55] = 32'h0;  // 32'hb86a3575;
    ram_cell[      56] = 32'h0;  // 32'h581e2d8f;
    ram_cell[      57] = 32'h0;  // 32'hdff6bd03;
    ram_cell[      58] = 32'h0;  // 32'h9926263e;
    ram_cell[      59] = 32'h0;  // 32'h7f8e7d9b;
    ram_cell[      60] = 32'h0;  // 32'h19378df1;
    ram_cell[      61] = 32'h0;  // 32'hd182a502;
    ram_cell[      62] = 32'h0;  // 32'h4ea3278d;
    ram_cell[      63] = 32'h0;  // 32'h8a31d7f6;
    ram_cell[      64] = 32'h0;  // 32'h37884312;
    ram_cell[      65] = 32'h0;  // 32'h15f65380;
    ram_cell[      66] = 32'h0;  // 32'h2ac9b80e;
    ram_cell[      67] = 32'h0;  // 32'h300f6b80;
    ram_cell[      68] = 32'h0;  // 32'h3530efa5;
    ram_cell[      69] = 32'h0;  // 32'hb4b15e10;
    ram_cell[      70] = 32'h0;  // 32'hecb014aa;
    ram_cell[      71] = 32'h0;  // 32'h178370a4;
    ram_cell[      72] = 32'h0;  // 32'h97bd6802;
    ram_cell[      73] = 32'h0;  // 32'h6e277ce1;
    ram_cell[      74] = 32'h0;  // 32'h5dd1d32a;
    ram_cell[      75] = 32'h0;  // 32'hf6da19b4;
    ram_cell[      76] = 32'h0;  // 32'hc34dbbb3;
    ram_cell[      77] = 32'h0;  // 32'hdd229ff1;
    ram_cell[      78] = 32'h0;  // 32'h6dd940cd;
    ram_cell[      79] = 32'h0;  // 32'h650809bd;
    ram_cell[      80] = 32'h0;  // 32'h5c9c1191;
    ram_cell[      81] = 32'h0;  // 32'h3e53c65b;
    ram_cell[      82] = 32'h0;  // 32'h0380c630;
    ram_cell[      83] = 32'h0;  // 32'h39a6ae0c;
    ram_cell[      84] = 32'h0;  // 32'h5ca59d69;
    ram_cell[      85] = 32'h0;  // 32'h7394045c;
    ram_cell[      86] = 32'h0;  // 32'h18b3483d;
    ram_cell[      87] = 32'h0;  // 32'h6a80fe58;
    ram_cell[      88] = 32'h0;  // 32'h8aa0f0e6;
    ram_cell[      89] = 32'h0;  // 32'hfd722db4;
    ram_cell[      90] = 32'h0;  // 32'h85082b9a;
    ram_cell[      91] = 32'h0;  // 32'hef05116f;
    ram_cell[      92] = 32'h0;  // 32'h68fbca8e;
    ram_cell[      93] = 32'h0;  // 32'h989924fd;
    ram_cell[      94] = 32'h0;  // 32'h06229382;
    ram_cell[      95] = 32'h0;  // 32'h4e94d0d6;
    ram_cell[      96] = 32'h0;  // 32'h0b6f34e0;
    ram_cell[      97] = 32'h0;  // 32'h3a1f8c66;
    ram_cell[      98] = 32'h0;  // 32'h9137cc06;
    ram_cell[      99] = 32'h0;  // 32'h87c81a6f;
    ram_cell[     100] = 32'h0;  // 32'h6acd896d;
    ram_cell[     101] = 32'h0;  // 32'hff827bc2;
    ram_cell[     102] = 32'h0;  // 32'hddacd22b;
    ram_cell[     103] = 32'h0;  // 32'hfbccbffb;
    ram_cell[     104] = 32'h0;  // 32'h3fe6bf79;
    ram_cell[     105] = 32'h0;  // 32'h3c967a4f;
    ram_cell[     106] = 32'h0;  // 32'h80b4fa4d;
    ram_cell[     107] = 32'h0;  // 32'h2cb462ae;
    ram_cell[     108] = 32'h0;  // 32'h58f3c0cd;
    ram_cell[     109] = 32'h0;  // 32'h9f345af8;
    ram_cell[     110] = 32'h0;  // 32'h7287aa31;
    ram_cell[     111] = 32'h0;  // 32'hc421656f;
    ram_cell[     112] = 32'h0;  // 32'hfb74d480;
    ram_cell[     113] = 32'h0;  // 32'h08ecedc1;
    ram_cell[     114] = 32'h0;  // 32'h5ef16c85;
    ram_cell[     115] = 32'h0;  // 32'h16789f5f;
    ram_cell[     116] = 32'h0;  // 32'hd59a5f11;
    ram_cell[     117] = 32'h0;  // 32'he687ca87;
    ram_cell[     118] = 32'h0;  // 32'hc63b0598;
    ram_cell[     119] = 32'h0;  // 32'h86244e13;
    ram_cell[     120] = 32'h0;  // 32'h52ae1070;
    ram_cell[     121] = 32'h0;  // 32'h6c1f33a7;
    ram_cell[     122] = 32'h0;  // 32'h0141ce8d;
    ram_cell[     123] = 32'h0;  // 32'h98e4e705;
    ram_cell[     124] = 32'h0;  // 32'h5587e6a4;
    ram_cell[     125] = 32'h0;  // 32'hbba97fae;
    ram_cell[     126] = 32'h0;  // 32'h0c26b2ab;
    ram_cell[     127] = 32'h0;  // 32'hc6502317;
    ram_cell[     128] = 32'h0;  // 32'h53a3aa98;
    ram_cell[     129] = 32'h0;  // 32'h6686500c;
    ram_cell[     130] = 32'h0;  // 32'h887a5b90;
    ram_cell[     131] = 32'h0;  // 32'h56e66662;
    ram_cell[     132] = 32'h0;  // 32'h67793beb;
    ram_cell[     133] = 32'h0;  // 32'h49e702d0;
    ram_cell[     134] = 32'h0;  // 32'h29ff0630;
    ram_cell[     135] = 32'h0;  // 32'hcdd1d6f0;
    ram_cell[     136] = 32'h0;  // 32'h1c726738;
    ram_cell[     137] = 32'h0;  // 32'h850d891f;
    ram_cell[     138] = 32'h0;  // 32'he0ae6822;
    ram_cell[     139] = 32'h0;  // 32'h998e35c9;
    ram_cell[     140] = 32'h0;  // 32'h4837b604;
    ram_cell[     141] = 32'h0;  // 32'h8c9d8d6c;
    ram_cell[     142] = 32'h0;  // 32'h8e2733b5;
    ram_cell[     143] = 32'h0;  // 32'ha026a8de;
    ram_cell[     144] = 32'h0;  // 32'hebacfd68;
    ram_cell[     145] = 32'h0;  // 32'h314a665f;
    ram_cell[     146] = 32'h0;  // 32'h18d99d95;
    ram_cell[     147] = 32'h0;  // 32'h5085eda7;
    ram_cell[     148] = 32'h0;  // 32'h7014baf9;
    ram_cell[     149] = 32'h0;  // 32'hc60b6450;
    ram_cell[     150] = 32'h0;  // 32'h60f0a445;
    ram_cell[     151] = 32'h0;  // 32'h20aae133;
    ram_cell[     152] = 32'h0;  // 32'h50ba1dcb;
    ram_cell[     153] = 32'h0;  // 32'h505cb7a5;
    ram_cell[     154] = 32'h0;  // 32'hd99e311b;
    ram_cell[     155] = 32'h0;  // 32'hfae8e162;
    ram_cell[     156] = 32'h0;  // 32'h67b0c60c;
    ram_cell[     157] = 32'h0;  // 32'hfd961459;
    ram_cell[     158] = 32'h0;  // 32'hc88a573b;
    ram_cell[     159] = 32'h0;  // 32'h7c89b746;
    ram_cell[     160] = 32'h0;  // 32'h6e7bfafc;
    ram_cell[     161] = 32'h0;  // 32'h4e12efbe;
    ram_cell[     162] = 32'h0;  // 32'h3709a6db;
    ram_cell[     163] = 32'h0;  // 32'h2d0b90c5;
    ram_cell[     164] = 32'h0;  // 32'he37ea8f2;
    ram_cell[     165] = 32'h0;  // 32'hd43e83f1;
    ram_cell[     166] = 32'h0;  // 32'h9600a44e;
    ram_cell[     167] = 32'h0;  // 32'hff133ac9;
    ram_cell[     168] = 32'h0;  // 32'h7f1f7821;
    ram_cell[     169] = 32'h0;  // 32'h77e9ee54;
    ram_cell[     170] = 32'h0;  // 32'h63d4fe81;
    ram_cell[     171] = 32'h0;  // 32'h5cbe74f8;
    ram_cell[     172] = 32'h0;  // 32'h2d347476;
    ram_cell[     173] = 32'h0;  // 32'h8bc8b52a;
    ram_cell[     174] = 32'h0;  // 32'hb19b987b;
    ram_cell[     175] = 32'h0;  // 32'hb8d60a68;
    ram_cell[     176] = 32'h0;  // 32'h4bea557f;
    ram_cell[     177] = 32'h0;  // 32'h8a437944;
    ram_cell[     178] = 32'h0;  // 32'h3bafbece;
    ram_cell[     179] = 32'h0;  // 32'h4abf4a3e;
    ram_cell[     180] = 32'h0;  // 32'h61cf2c51;
    ram_cell[     181] = 32'h0;  // 32'h6db0982d;
    ram_cell[     182] = 32'h0;  // 32'h6863eb52;
    ram_cell[     183] = 32'h0;  // 32'h03086bc0;
    ram_cell[     184] = 32'h0;  // 32'hb277234a;
    ram_cell[     185] = 32'h0;  // 32'h0eee9561;
    ram_cell[     186] = 32'h0;  // 32'h0b747bef;
    ram_cell[     187] = 32'h0;  // 32'hba0600ed;
    ram_cell[     188] = 32'h0;  // 32'h78d39140;
    ram_cell[     189] = 32'h0;  // 32'hfcce770f;
    ram_cell[     190] = 32'h0;  // 32'h36c36423;
    ram_cell[     191] = 32'h0;  // 32'h15f46818;
    ram_cell[     192] = 32'h0;  // 32'h9543eb27;
    ram_cell[     193] = 32'h0;  // 32'hcce63efd;
    ram_cell[     194] = 32'h0;  // 32'h5304d48c;
    ram_cell[     195] = 32'h0;  // 32'h1649b3a6;
    ram_cell[     196] = 32'h0;  // 32'hfb8562a6;
    ram_cell[     197] = 32'h0;  // 32'h840e1eef;
    ram_cell[     198] = 32'h0;  // 32'hbac135b6;
    ram_cell[     199] = 32'h0;  // 32'h26027469;
    ram_cell[     200] = 32'h0;  // 32'h3d90b349;
    ram_cell[     201] = 32'h0;  // 32'h6631467c;
    ram_cell[     202] = 32'h0;  // 32'ha0b3fb63;
    ram_cell[     203] = 32'h0;  // 32'h10cb9582;
    ram_cell[     204] = 32'h0;  // 32'h6c43b7c2;
    ram_cell[     205] = 32'h0;  // 32'h10fb1cef;
    ram_cell[     206] = 32'h0;  // 32'h12237a4d;
    ram_cell[     207] = 32'h0;  // 32'h33051968;
    ram_cell[     208] = 32'h0;  // 32'h2b214b18;
    ram_cell[     209] = 32'h0;  // 32'h9f385d25;
    ram_cell[     210] = 32'h0;  // 32'h49f24282;
    ram_cell[     211] = 32'h0;  // 32'h5a927dc8;
    ram_cell[     212] = 32'h0;  // 32'h153125ef;
    ram_cell[     213] = 32'h0;  // 32'h08cb9a2f;
    ram_cell[     214] = 32'h0;  // 32'hca7f6560;
    ram_cell[     215] = 32'h0;  // 32'h9fe0af67;
    ram_cell[     216] = 32'h0;  // 32'ha55fe45d;
    ram_cell[     217] = 32'h0;  // 32'h495fffaf;
    ram_cell[     218] = 32'h0;  // 32'h92e43c7c;
    ram_cell[     219] = 32'h0;  // 32'h22a0de5c;
    ram_cell[     220] = 32'h0;  // 32'h5421949e;
    ram_cell[     221] = 32'h0;  // 32'had042ae1;
    ram_cell[     222] = 32'h0;  // 32'h5e99121b;
    ram_cell[     223] = 32'h0;  // 32'hb1917fe7;
    ram_cell[     224] = 32'h0;  // 32'h57708f53;
    ram_cell[     225] = 32'h0;  // 32'h3d4d4744;
    ram_cell[     226] = 32'h0;  // 32'h4408ccbd;
    ram_cell[     227] = 32'h0;  // 32'h423312b3;
    ram_cell[     228] = 32'h0;  // 32'hbf439e56;
    ram_cell[     229] = 32'h0;  // 32'h7d7d5781;
    ram_cell[     230] = 32'h0;  // 32'h2666c916;
    ram_cell[     231] = 32'h0;  // 32'hfff0edcd;
    ram_cell[     232] = 32'h0;  // 32'h40235176;
    ram_cell[     233] = 32'h0;  // 32'h8e2852d2;
    ram_cell[     234] = 32'h0;  // 32'h49efb7d2;
    ram_cell[     235] = 32'h0;  // 32'ha78c9ccf;
    ram_cell[     236] = 32'h0;  // 32'h7e170600;
    ram_cell[     237] = 32'h0;  // 32'h0dda948d;
    ram_cell[     238] = 32'h0;  // 32'h7df7bdea;
    ram_cell[     239] = 32'h0;  // 32'h81f318d7;
    ram_cell[     240] = 32'h0;  // 32'hd1d4d9fe;
    ram_cell[     241] = 32'h0;  // 32'h458a8f0f;
    ram_cell[     242] = 32'h0;  // 32'hc794d7b0;
    ram_cell[     243] = 32'h0;  // 32'hcf9c9f00;
    ram_cell[     244] = 32'h0;  // 32'h870bd653;
    ram_cell[     245] = 32'h0;  // 32'h6d6cdcdf;
    ram_cell[     246] = 32'h0;  // 32'h303fdb0d;
    ram_cell[     247] = 32'h0;  // 32'h9b7fd19c;
    ram_cell[     248] = 32'h0;  // 32'hd421bdae;
    ram_cell[     249] = 32'h0;  // 32'hc005cb45;
    ram_cell[     250] = 32'h0;  // 32'h399a3704;
    ram_cell[     251] = 32'h0;  // 32'hec648090;
    ram_cell[     252] = 32'h0;  // 32'ha9dc7a34;
    ram_cell[     253] = 32'h0;  // 32'h9c506a6e;
    ram_cell[     254] = 32'h0;  // 32'h08c7883b;
    ram_cell[     255] = 32'h0;  // 32'h46a5bbac;
    // src matrix A
    ram_cell[     256] = 32'hbcef2b9b;
    ram_cell[     257] = 32'ha88f34cd;
    ram_cell[     258] = 32'h37b33170;
    ram_cell[     259] = 32'hae74868b;
    ram_cell[     260] = 32'h97cbf93d;
    ram_cell[     261] = 32'hb2988fa8;
    ram_cell[     262] = 32'hb23970ac;
    ram_cell[     263] = 32'h6ace8384;
    ram_cell[     264] = 32'h7af5d5c7;
    ram_cell[     265] = 32'h29c40856;
    ram_cell[     266] = 32'ha2d817e1;
    ram_cell[     267] = 32'hc49040ce;
    ram_cell[     268] = 32'hf7664d20;
    ram_cell[     269] = 32'hdbd52faa;
    ram_cell[     270] = 32'h4e07cfd4;
    ram_cell[     271] = 32'hf031f510;
    ram_cell[     272] = 32'hf444358c;
    ram_cell[     273] = 32'hda326c13;
    ram_cell[     274] = 32'h701d1338;
    ram_cell[     275] = 32'h6b5d65d9;
    ram_cell[     276] = 32'had2e5d5a;
    ram_cell[     277] = 32'h34286eea;
    ram_cell[     278] = 32'h461cfcb2;
    ram_cell[     279] = 32'hf3682cfe;
    ram_cell[     280] = 32'h60a7cada;
    ram_cell[     281] = 32'h8b742378;
    ram_cell[     282] = 32'h2ac7cf2c;
    ram_cell[     283] = 32'h32d0d124;
    ram_cell[     284] = 32'h5d80e631;
    ram_cell[     285] = 32'h667b47ce;
    ram_cell[     286] = 32'ha97d5c38;
    ram_cell[     287] = 32'h7343c12e;
    ram_cell[     288] = 32'h3c3129d6;
    ram_cell[     289] = 32'h6cdb5ef3;
    ram_cell[     290] = 32'h2194df1a;
    ram_cell[     291] = 32'h117b5b08;
    ram_cell[     292] = 32'h9de589d1;
    ram_cell[     293] = 32'h0451d5f1;
    ram_cell[     294] = 32'heb7b843a;
    ram_cell[     295] = 32'he643c1e0;
    ram_cell[     296] = 32'hacbd54ff;
    ram_cell[     297] = 32'hab20b829;
    ram_cell[     298] = 32'hc01a541f;
    ram_cell[     299] = 32'ha9234053;
    ram_cell[     300] = 32'h90e544f8;
    ram_cell[     301] = 32'h6b1eb2fe;
    ram_cell[     302] = 32'h3a507d58;
    ram_cell[     303] = 32'h0f53d721;
    ram_cell[     304] = 32'h0125ee87;
    ram_cell[     305] = 32'h9c4e2d7d;
    ram_cell[     306] = 32'hb9e20050;
    ram_cell[     307] = 32'h044a9bc0;
    ram_cell[     308] = 32'h6b396da7;
    ram_cell[     309] = 32'h32701891;
    ram_cell[     310] = 32'h372bde57;
    ram_cell[     311] = 32'h3654b666;
    ram_cell[     312] = 32'h5aa200c5;
    ram_cell[     313] = 32'hc5413f83;
    ram_cell[     314] = 32'h956623b3;
    ram_cell[     315] = 32'hf631a2c4;
    ram_cell[     316] = 32'hfced0025;
    ram_cell[     317] = 32'h795be146;
    ram_cell[     318] = 32'he427e332;
    ram_cell[     319] = 32'hbb8013bf;
    ram_cell[     320] = 32'h33a40750;
    ram_cell[     321] = 32'h4a73a541;
    ram_cell[     322] = 32'h45374da8;
    ram_cell[     323] = 32'hdf71ccc5;
    ram_cell[     324] = 32'h11a75dd3;
    ram_cell[     325] = 32'h7c8db6d9;
    ram_cell[     326] = 32'h28396b2e;
    ram_cell[     327] = 32'h2d9012c3;
    ram_cell[     328] = 32'hfc790691;
    ram_cell[     329] = 32'he8e0e287;
    ram_cell[     330] = 32'h4a360b44;
    ram_cell[     331] = 32'hb7bedbe1;
    ram_cell[     332] = 32'h7f12691a;
    ram_cell[     333] = 32'h8a9c515b;
    ram_cell[     334] = 32'h5ac41e5e;
    ram_cell[     335] = 32'h9318ec9a;
    ram_cell[     336] = 32'h15dfd15c;
    ram_cell[     337] = 32'h4e7feaf2;
    ram_cell[     338] = 32'hea95346d;
    ram_cell[     339] = 32'hbda29a15;
    ram_cell[     340] = 32'h514ce4ad;
    ram_cell[     341] = 32'h0679f706;
    ram_cell[     342] = 32'h1fef36ea;
    ram_cell[     343] = 32'h857b5e3b;
    ram_cell[     344] = 32'h7bbd9726;
    ram_cell[     345] = 32'haeda0bd1;
    ram_cell[     346] = 32'h4d6c474b;
    ram_cell[     347] = 32'ha16761cc;
    ram_cell[     348] = 32'h29fe3231;
    ram_cell[     349] = 32'h3ab4aaf4;
    ram_cell[     350] = 32'h9f5d36e2;
    ram_cell[     351] = 32'hc53e46b3;
    ram_cell[     352] = 32'h25b2cc79;
    ram_cell[     353] = 32'h2c113e27;
    ram_cell[     354] = 32'h13196927;
    ram_cell[     355] = 32'h2d78ca04;
    ram_cell[     356] = 32'h861f397c;
    ram_cell[     357] = 32'h164db1e4;
    ram_cell[     358] = 32'h786a324a;
    ram_cell[     359] = 32'he28ed383;
    ram_cell[     360] = 32'ha55f1615;
    ram_cell[     361] = 32'hb892298b;
    ram_cell[     362] = 32'hb35f662b;
    ram_cell[     363] = 32'hd6155bb4;
    ram_cell[     364] = 32'h9f8e9e72;
    ram_cell[     365] = 32'h78185039;
    ram_cell[     366] = 32'h69d9d649;
    ram_cell[     367] = 32'h4595faed;
    ram_cell[     368] = 32'h862a3263;
    ram_cell[     369] = 32'h6d504d69;
    ram_cell[     370] = 32'h211df87b;
    ram_cell[     371] = 32'h1c588ffd;
    ram_cell[     372] = 32'h1c4a796b;
    ram_cell[     373] = 32'h94ea41e2;
    ram_cell[     374] = 32'h10c24992;
    ram_cell[     375] = 32'hb8b8818e;
    ram_cell[     376] = 32'h71867513;
    ram_cell[     377] = 32'h292ddb0a;
    ram_cell[     378] = 32'he1d7d03f;
    ram_cell[     379] = 32'hb60d5727;
    ram_cell[     380] = 32'h41e00a03;
    ram_cell[     381] = 32'h55c28962;
    ram_cell[     382] = 32'h2e42208f;
    ram_cell[     383] = 32'h8b27a81b;
    ram_cell[     384] = 32'h4e470d34;
    ram_cell[     385] = 32'h4beecd41;
    ram_cell[     386] = 32'h34e33d4b;
    ram_cell[     387] = 32'he83580a4;
    ram_cell[     388] = 32'h43cd04c5;
    ram_cell[     389] = 32'h3d194c23;
    ram_cell[     390] = 32'heb4097a9;
    ram_cell[     391] = 32'h343ee732;
    ram_cell[     392] = 32'h33af291f;
    ram_cell[     393] = 32'h96f519a1;
    ram_cell[     394] = 32'h0d924ff9;
    ram_cell[     395] = 32'h2ff0e755;
    ram_cell[     396] = 32'hb52c7839;
    ram_cell[     397] = 32'h792ad159;
    ram_cell[     398] = 32'h4e2d64eb;
    ram_cell[     399] = 32'he70a795c;
    ram_cell[     400] = 32'h7e8bfe19;
    ram_cell[     401] = 32'h2ceaf97b;
    ram_cell[     402] = 32'h6c1e5016;
    ram_cell[     403] = 32'hc6c96042;
    ram_cell[     404] = 32'h1d024f00;
    ram_cell[     405] = 32'h467546a7;
    ram_cell[     406] = 32'ha44a93c3;
    ram_cell[     407] = 32'h126c853c;
    ram_cell[     408] = 32'hb8ce9041;
    ram_cell[     409] = 32'h7876f057;
    ram_cell[     410] = 32'h65fa7da8;
    ram_cell[     411] = 32'hbe245dbe;
    ram_cell[     412] = 32'h2ab9d9b3;
    ram_cell[     413] = 32'h79e4153b;
    ram_cell[     414] = 32'h8fcd66d8;
    ram_cell[     415] = 32'h57f36967;
    ram_cell[     416] = 32'h1c8baf9a;
    ram_cell[     417] = 32'h03b896a0;
    ram_cell[     418] = 32'h85f7aec7;
    ram_cell[     419] = 32'hc8b5650f;
    ram_cell[     420] = 32'h09b77cdb;
    ram_cell[     421] = 32'h2318047e;
    ram_cell[     422] = 32'h1de6d34a;
    ram_cell[     423] = 32'he56e915c;
    ram_cell[     424] = 32'hf93e5170;
    ram_cell[     425] = 32'h8d1ede91;
    ram_cell[     426] = 32'hf03f8dec;
    ram_cell[     427] = 32'h0df757b0;
    ram_cell[     428] = 32'hb5a38e66;
    ram_cell[     429] = 32'he8718af0;
    ram_cell[     430] = 32'h793bcf1b;
    ram_cell[     431] = 32'hac4cbec0;
    ram_cell[     432] = 32'h752b0f05;
    ram_cell[     433] = 32'h46d3d286;
    ram_cell[     434] = 32'hb19ed556;
    ram_cell[     435] = 32'ha04aca3d;
    ram_cell[     436] = 32'h625556a3;
    ram_cell[     437] = 32'hfbf320fe;
    ram_cell[     438] = 32'h4d75bdab;
    ram_cell[     439] = 32'h7d412065;
    ram_cell[     440] = 32'h9e1c5294;
    ram_cell[     441] = 32'h26c681da;
    ram_cell[     442] = 32'hb17b4a78;
    ram_cell[     443] = 32'ha8f3d641;
    ram_cell[     444] = 32'ha742d5e5;
    ram_cell[     445] = 32'heee5029a;
    ram_cell[     446] = 32'h43f93b7f;
    ram_cell[     447] = 32'h515937c9;
    ram_cell[     448] = 32'h44cb2435;
    ram_cell[     449] = 32'hcb1e9c87;
    ram_cell[     450] = 32'h3bf116c7;
    ram_cell[     451] = 32'he5037812;
    ram_cell[     452] = 32'h4be05f91;
    ram_cell[     453] = 32'h14cd0ac2;
    ram_cell[     454] = 32'h2054953e;
    ram_cell[     455] = 32'h710bacfb;
    ram_cell[     456] = 32'haf1b2725;
    ram_cell[     457] = 32'h53574fa4;
    ram_cell[     458] = 32'hab9d5c5f;
    ram_cell[     459] = 32'h9f0731ef;
    ram_cell[     460] = 32'hf86fdf52;
    ram_cell[     461] = 32'he7d81a44;
    ram_cell[     462] = 32'h558aca30;
    ram_cell[     463] = 32'h826a79fa;
    ram_cell[     464] = 32'h0c54820d;
    ram_cell[     465] = 32'hc5318ff6;
    ram_cell[     466] = 32'h83c5a55a;
    ram_cell[     467] = 32'h43150486;
    ram_cell[     468] = 32'h0ce7c1d9;
    ram_cell[     469] = 32'he7232ee0;
    ram_cell[     470] = 32'h61825999;
    ram_cell[     471] = 32'hb3c8b614;
    ram_cell[     472] = 32'h5d2572cd;
    ram_cell[     473] = 32'h473e7c28;
    ram_cell[     474] = 32'h73338da5;
    ram_cell[     475] = 32'h64d3e5ff;
    ram_cell[     476] = 32'hc53981ae;
    ram_cell[     477] = 32'hd8bec2f2;
    ram_cell[     478] = 32'h78e1e4e4;
    ram_cell[     479] = 32'hca50fe66;
    ram_cell[     480] = 32'h46a76928;
    ram_cell[     481] = 32'h41249954;
    ram_cell[     482] = 32'he73edcec;
    ram_cell[     483] = 32'hec42ffc3;
    ram_cell[     484] = 32'hb33d4718;
    ram_cell[     485] = 32'hba421df1;
    ram_cell[     486] = 32'hf8ecdf10;
    ram_cell[     487] = 32'h60aeeba4;
    ram_cell[     488] = 32'hbfa0aeaa;
    ram_cell[     489] = 32'hd43a2049;
    ram_cell[     490] = 32'h172447b9;
    ram_cell[     491] = 32'he44af5b7;
    ram_cell[     492] = 32'h69380693;
    ram_cell[     493] = 32'h321e4db2;
    ram_cell[     494] = 32'hd32d0034;
    ram_cell[     495] = 32'hc6802feb;
    ram_cell[     496] = 32'h5e3b8fe4;
    ram_cell[     497] = 32'h5d2d6871;
    ram_cell[     498] = 32'h1fa4e4cf;
    ram_cell[     499] = 32'h25cfd8b8;
    ram_cell[     500] = 32'h3ff71ac5;
    ram_cell[     501] = 32'h625c0b35;
    ram_cell[     502] = 32'ha26dbea1;
    ram_cell[     503] = 32'h5d87c2cd;
    ram_cell[     504] = 32'hdb1407f4;
    ram_cell[     505] = 32'heb762597;
    ram_cell[     506] = 32'h23540f63;
    ram_cell[     507] = 32'hac619fdf;
    ram_cell[     508] = 32'h442e7a33;
    ram_cell[     509] = 32'h52d49971;
    ram_cell[     510] = 32'h67c4e1e8;
    ram_cell[     511] = 32'h504edaa4;
    // src matrix B
    ram_cell[     512] = 32'h8366e20c;
    ram_cell[     513] = 32'h77659227;
    ram_cell[     514] = 32'h2599174a;
    ram_cell[     515] = 32'h91b7973c;
    ram_cell[     516] = 32'h14e1a28d;
    ram_cell[     517] = 32'h38bd5572;
    ram_cell[     518] = 32'h6f5ea0de;
    ram_cell[     519] = 32'h0d2b0c75;
    ram_cell[     520] = 32'h0b1e6396;
    ram_cell[     521] = 32'h17f6c35f;
    ram_cell[     522] = 32'h4f801e52;
    ram_cell[     523] = 32'hce4f651c;
    ram_cell[     524] = 32'hcbf2fe27;
    ram_cell[     525] = 32'ha3dd0d4b;
    ram_cell[     526] = 32'hf91fe10b;
    ram_cell[     527] = 32'ha092f6c4;
    ram_cell[     528] = 32'h3158fd79;
    ram_cell[     529] = 32'h1a1ce404;
    ram_cell[     530] = 32'hac57bead;
    ram_cell[     531] = 32'h8770e0f3;
    ram_cell[     532] = 32'h4d876912;
    ram_cell[     533] = 32'h73dfa643;
    ram_cell[     534] = 32'h2cdf14d5;
    ram_cell[     535] = 32'ha5617030;
    ram_cell[     536] = 32'hf986f114;
    ram_cell[     537] = 32'h238e674b;
    ram_cell[     538] = 32'he9c94e57;
    ram_cell[     539] = 32'hf02cd770;
    ram_cell[     540] = 32'hf649ae25;
    ram_cell[     541] = 32'h686c55e8;
    ram_cell[     542] = 32'he644dabf;
    ram_cell[     543] = 32'h909e749b;
    ram_cell[     544] = 32'h4081d82c;
    ram_cell[     545] = 32'h774113ab;
    ram_cell[     546] = 32'h69db6e16;
    ram_cell[     547] = 32'h9a856630;
    ram_cell[     548] = 32'h3e4ae39b;
    ram_cell[     549] = 32'h8dc098ca;
    ram_cell[     550] = 32'h5a683173;
    ram_cell[     551] = 32'h0b21bf21;
    ram_cell[     552] = 32'hf9ef5fb4;
    ram_cell[     553] = 32'hc840c965;
    ram_cell[     554] = 32'h8940bcc0;
    ram_cell[     555] = 32'hcaffc505;
    ram_cell[     556] = 32'h81a597bd;
    ram_cell[     557] = 32'hddbecddd;
    ram_cell[     558] = 32'h4c453bd9;
    ram_cell[     559] = 32'hdd53cc6e;
    ram_cell[     560] = 32'hc7263e04;
    ram_cell[     561] = 32'he6e283b3;
    ram_cell[     562] = 32'h7a935c98;
    ram_cell[     563] = 32'hc987bb37;
    ram_cell[     564] = 32'h7ef4f00d;
    ram_cell[     565] = 32'h32b41671;
    ram_cell[     566] = 32'h60d3be00;
    ram_cell[     567] = 32'he18e5912;
    ram_cell[     568] = 32'h4177262d;
    ram_cell[     569] = 32'hc9da93ef;
    ram_cell[     570] = 32'h1e8d59a3;
    ram_cell[     571] = 32'ha727c825;
    ram_cell[     572] = 32'h0f9e659a;
    ram_cell[     573] = 32'h16c1c661;
    ram_cell[     574] = 32'h1b8ccbc3;
    ram_cell[     575] = 32'h4c939ce4;
    ram_cell[     576] = 32'hb9cc7b0e;
    ram_cell[     577] = 32'he0eeadf8;
    ram_cell[     578] = 32'h9850aa4c;
    ram_cell[     579] = 32'hd0d8bdb8;
    ram_cell[     580] = 32'hd383a3df;
    ram_cell[     581] = 32'hc2108b2b;
    ram_cell[     582] = 32'h29e06220;
    ram_cell[     583] = 32'he3952675;
    ram_cell[     584] = 32'hb2a47d1b;
    ram_cell[     585] = 32'h116d4672;
    ram_cell[     586] = 32'hac017848;
    ram_cell[     587] = 32'h50c3e653;
    ram_cell[     588] = 32'h5dc7b8a6;
    ram_cell[     589] = 32'h0edfffb7;
    ram_cell[     590] = 32'hd43c9e5c;
    ram_cell[     591] = 32'h8abb2ed2;
    ram_cell[     592] = 32'hb28abfea;
    ram_cell[     593] = 32'hfaa037f2;
    ram_cell[     594] = 32'h633753e3;
    ram_cell[     595] = 32'h525b6519;
    ram_cell[     596] = 32'h17856329;
    ram_cell[     597] = 32'he94d8b0f;
    ram_cell[     598] = 32'h89ec497c;
    ram_cell[     599] = 32'h16c59466;
    ram_cell[     600] = 32'h91d8646d;
    ram_cell[     601] = 32'hfe6ccf45;
    ram_cell[     602] = 32'h5ff99615;
    ram_cell[     603] = 32'h7ac22270;
    ram_cell[     604] = 32'h89315e2e;
    ram_cell[     605] = 32'h07c27f25;
    ram_cell[     606] = 32'h21fbb6ad;
    ram_cell[     607] = 32'hd4521714;
    ram_cell[     608] = 32'h661a3b7b;
    ram_cell[     609] = 32'hb7daf3d4;
    ram_cell[     610] = 32'ha9ba0eed;
    ram_cell[     611] = 32'hfaa4c172;
    ram_cell[     612] = 32'hb3b26a3f;
    ram_cell[     613] = 32'h13641785;
    ram_cell[     614] = 32'h91bf0361;
    ram_cell[     615] = 32'hb7f98302;
    ram_cell[     616] = 32'he3cb2dfc;
    ram_cell[     617] = 32'hb2cb8f51;
    ram_cell[     618] = 32'h221fbcdd;
    ram_cell[     619] = 32'ha8c11962;
    ram_cell[     620] = 32'h15f03bfb;
    ram_cell[     621] = 32'h7c801b1a;
    ram_cell[     622] = 32'hee3e4601;
    ram_cell[     623] = 32'h83f546ec;
    ram_cell[     624] = 32'hf0eecebb;
    ram_cell[     625] = 32'h26e6de39;
    ram_cell[     626] = 32'hda620104;
    ram_cell[     627] = 32'h451af5d9;
    ram_cell[     628] = 32'h780d0f0f;
    ram_cell[     629] = 32'h92887d60;
    ram_cell[     630] = 32'h268c4e51;
    ram_cell[     631] = 32'he109b0c3;
    ram_cell[     632] = 32'h8763a43e;
    ram_cell[     633] = 32'hb61837b6;
    ram_cell[     634] = 32'h6bfced43;
    ram_cell[     635] = 32'h5c3a8e6b;
    ram_cell[     636] = 32'h73276d65;
    ram_cell[     637] = 32'ha05a981b;
    ram_cell[     638] = 32'he3690f4b;
    ram_cell[     639] = 32'h8533ed08;
    ram_cell[     640] = 32'hd87f49fa;
    ram_cell[     641] = 32'hdfb540f1;
    ram_cell[     642] = 32'h7c3705df;
    ram_cell[     643] = 32'he453eb2a;
    ram_cell[     644] = 32'h4afe9900;
    ram_cell[     645] = 32'h71035e94;
    ram_cell[     646] = 32'hc79c0bb5;
    ram_cell[     647] = 32'h03c1fa28;
    ram_cell[     648] = 32'h56196b19;
    ram_cell[     649] = 32'h8b4dfcf1;
    ram_cell[     650] = 32'h2522a9ab;
    ram_cell[     651] = 32'hbd0edd01;
    ram_cell[     652] = 32'h12130c36;
    ram_cell[     653] = 32'hca1f27c8;
    ram_cell[     654] = 32'h03d18dc4;
    ram_cell[     655] = 32'h25d2f9df;
    ram_cell[     656] = 32'h7cd044e3;
    ram_cell[     657] = 32'h9dd89def;
    ram_cell[     658] = 32'hfb3dbeb2;
    ram_cell[     659] = 32'h0c33a0a5;
    ram_cell[     660] = 32'h0c61e626;
    ram_cell[     661] = 32'h690b9264;
    ram_cell[     662] = 32'ha2fdcd18;
    ram_cell[     663] = 32'h530ae0c2;
    ram_cell[     664] = 32'h0e96961e;
    ram_cell[     665] = 32'h0789f69b;
    ram_cell[     666] = 32'hb4a081be;
    ram_cell[     667] = 32'h3d91e1e6;
    ram_cell[     668] = 32'h4dd04a1e;
    ram_cell[     669] = 32'h944337ea;
    ram_cell[     670] = 32'h28fbaf42;
    ram_cell[     671] = 32'hbbe2f819;
    ram_cell[     672] = 32'hb2195312;
    ram_cell[     673] = 32'h2a14def6;
    ram_cell[     674] = 32'hde2b3c7e;
    ram_cell[     675] = 32'hffc911bf;
    ram_cell[     676] = 32'h73c0ade3;
    ram_cell[     677] = 32'h8e94ac54;
    ram_cell[     678] = 32'h7ffd789d;
    ram_cell[     679] = 32'h885b5b2d;
    ram_cell[     680] = 32'hc0ae4895;
    ram_cell[     681] = 32'hf29707aa;
    ram_cell[     682] = 32'hc1c3c5fa;
    ram_cell[     683] = 32'h800c8f13;
    ram_cell[     684] = 32'h40943226;
    ram_cell[     685] = 32'hd4185219;
    ram_cell[     686] = 32'h8de2ad6e;
    ram_cell[     687] = 32'hdd74e501;
    ram_cell[     688] = 32'hfd0891e9;
    ram_cell[     689] = 32'hc7e8eca1;
    ram_cell[     690] = 32'hb66f06ee;
    ram_cell[     691] = 32'h53081801;
    ram_cell[     692] = 32'hbee5a3eb;
    ram_cell[     693] = 32'ha1e7d169;
    ram_cell[     694] = 32'hc968db17;
    ram_cell[     695] = 32'hd5b889ca;
    ram_cell[     696] = 32'h0a5e6e56;
    ram_cell[     697] = 32'h2da9adb4;
    ram_cell[     698] = 32'h5fbebfde;
    ram_cell[     699] = 32'h650c268b;
    ram_cell[     700] = 32'h873e0f3e;
    ram_cell[     701] = 32'h0fa1fe82;
    ram_cell[     702] = 32'hd024ba91;
    ram_cell[     703] = 32'hcd70eb11;
    ram_cell[     704] = 32'h55d3f83d;
    ram_cell[     705] = 32'hb6d24c74;
    ram_cell[     706] = 32'hf0b6f098;
    ram_cell[     707] = 32'h7965f3dc;
    ram_cell[     708] = 32'he85cf348;
    ram_cell[     709] = 32'h338f6e77;
    ram_cell[     710] = 32'hc4905b8f;
    ram_cell[     711] = 32'h02cdc1a0;
    ram_cell[     712] = 32'h7f13c307;
    ram_cell[     713] = 32'hd9ad7498;
    ram_cell[     714] = 32'hdc0f8e89;
    ram_cell[     715] = 32'h145617b8;
    ram_cell[     716] = 32'hfe4bbe21;
    ram_cell[     717] = 32'h6b659870;
    ram_cell[     718] = 32'hc961471d;
    ram_cell[     719] = 32'h3ae7b4ad;
    ram_cell[     720] = 32'hf46c6e0e;
    ram_cell[     721] = 32'h9389d76f;
    ram_cell[     722] = 32'h6c519ecb;
    ram_cell[     723] = 32'hb460036c;
    ram_cell[     724] = 32'h302d8e88;
    ram_cell[     725] = 32'ha4fcc5af;
    ram_cell[     726] = 32'hc47c26c4;
    ram_cell[     727] = 32'h728086e2;
    ram_cell[     728] = 32'h67fc185e;
    ram_cell[     729] = 32'h8bbf3c24;
    ram_cell[     730] = 32'h66200eef;
    ram_cell[     731] = 32'h505d7933;
    ram_cell[     732] = 32'he18ed0d1;
    ram_cell[     733] = 32'h09fcf331;
    ram_cell[     734] = 32'hd7d8024c;
    ram_cell[     735] = 32'h26c1b091;
    ram_cell[     736] = 32'h5fee4021;
    ram_cell[     737] = 32'h507aa05b;
    ram_cell[     738] = 32'hf8ca8125;
    ram_cell[     739] = 32'h27c2620b;
    ram_cell[     740] = 32'hf9421e65;
    ram_cell[     741] = 32'h8ba37709;
    ram_cell[     742] = 32'h8e8803e7;
    ram_cell[     743] = 32'h2f2b67d5;
    ram_cell[     744] = 32'hd06c54ad;
    ram_cell[     745] = 32'h9df33e03;
    ram_cell[     746] = 32'hd6729684;
    ram_cell[     747] = 32'h24b8e0bd;
    ram_cell[     748] = 32'h20dd0323;
    ram_cell[     749] = 32'h670a36ed;
    ram_cell[     750] = 32'h17814361;
    ram_cell[     751] = 32'h856d64c7;
    ram_cell[     752] = 32'hae799f78;
    ram_cell[     753] = 32'h14599545;
    ram_cell[     754] = 32'hdc952da2;
    ram_cell[     755] = 32'ha04655ca;
    ram_cell[     756] = 32'h02ac5d94;
    ram_cell[     757] = 32'ha806eb49;
    ram_cell[     758] = 32'h53464e7b;
    ram_cell[     759] = 32'h34d08e42;
    ram_cell[     760] = 32'h73db9d24;
    ram_cell[     761] = 32'hd1c6b3a9;
    ram_cell[     762] = 32'he87930ff;
    ram_cell[     763] = 32'h72e6cd08;
    ram_cell[     764] = 32'h1368a129;
    ram_cell[     765] = 32'h8bab6138;
    ram_cell[     766] = 32'ha23a5be4;
    ram_cell[     767] = 32'h82d5d1d5;
end

endmodule

