`timescale 1ns/100ps
//correct read result:
// 00000000 000000ef 00000048 00000129 000000e3 0000012e 00000135 00000008 000000a4 00000068 00000006 00000075 00000147 000000a7 00000188 0000011e 000000e9 0000009d 00000065 00000087 00000119 0000002e 00000010 000000fe 00000057 00000161 0000008a 000000ba 0000002e 000000a3 00000115 00000127 0000016e 000000f9 0000001c 00000059 00000067 0000011e 00000036 00000098 0000005f 0000015d 000000c1 0000014d 00000134 000000ff 00000136 00000173 0000007f 0000003e 0000001e 00000144 000000b0 0000014d 00000111 00000027 000000f9 00000123 00000163 00000046 0000002f 0000013f 000000ad 0000001d 0000015e 00000146 00000054 000000b0 0000015e 000000fa 00000173 0000008b 0000005d 00000117 0000015f 000000aa 00000156 00000138 00000000 000000f4 00000142 000000d5 000000ba 00000056 000000f9 000000ef 00000022 00000021 00000013 000000bf 00000091 000000e1 0000014d 0000001b 00000085 000000ad 000000c1 00000171 0000005d 00000009

module cache_tb();

`define DATA_COUNT (100)
`define RDWR_COUNT (6*`DATA_COUNT)

reg wr_cycle           [`RDWR_COUNT];
reg rd_cycle           [`RDWR_COUNT];
reg [31:0] addr_rom    [`RDWR_COUNT];
reg [31:0] wr_data_rom [`RDWR_COUNT];
reg [31:0] validation_data [`DATA_COUNT];

initial begin
    // 100 sequence write cycles
    rd_cycle[    0] = 1'b0;  wr_cycle[    0] = 1'b1;  addr_rom[    0]='h00000000;  wr_data_rom[    0]='h00000000;
    rd_cycle[    1] = 1'b0;  wr_cycle[    1] = 1'b1;  addr_rom[    1]='h00000004;  wr_data_rom[    1]='h0000005a;
    rd_cycle[    2] = 1'b0;  wr_cycle[    2] = 1'b1;  addr_rom[    2]='h00000008;  wr_data_rom[    2]='h00000048;
    rd_cycle[    3] = 1'b0;  wr_cycle[    3] = 1'b1;  addr_rom[    3]='h0000000c;  wr_data_rom[    3]='h000000fd;
    rd_cycle[    4] = 1'b0;  wr_cycle[    4] = 1'b1;  addr_rom[    4]='h00000010;  wr_data_rom[    4]='h000000e3;
    rd_cycle[    5] = 1'b0;  wr_cycle[    5] = 1'b1;  addr_rom[    5]='h00000014;  wr_data_rom[    5]='h0000012e;
    rd_cycle[    6] = 1'b0;  wr_cycle[    6] = 1'b1;  addr_rom[    6]='h00000018;  wr_data_rom[    6]='h00000178;
    rd_cycle[    7] = 1'b0;  wr_cycle[    7] = 1'b1;  addr_rom[    7]='h0000001c;  wr_data_rom[    7]='h0000011c;
    rd_cycle[    8] = 1'b0;  wr_cycle[    8] = 1'b1;  addr_rom[    8]='h00000020;  wr_data_rom[    8]='h00000124;
    rd_cycle[    9] = 1'b0;  wr_cycle[    9] = 1'b1;  addr_rom[    9]='h00000024;  wr_data_rom[    9]='h0000010b;
    rd_cycle[   10] = 1'b0;  wr_cycle[   10] = 1'b1;  addr_rom[   10]='h00000028;  wr_data_rom[   10]='h0000015a;
    rd_cycle[   11] = 1'b0;  wr_cycle[   11] = 1'b1;  addr_rom[   11]='h0000002c;  wr_data_rom[   11]='h00000189;
    rd_cycle[   12] = 1'b0;  wr_cycle[   12] = 1'b1;  addr_rom[   12]='h00000030;  wr_data_rom[   12]='h00000052;
    rd_cycle[   13] = 1'b0;  wr_cycle[   13] = 1'b1;  addr_rom[   13]='h00000034;  wr_data_rom[   13]='h000000a7;
    rd_cycle[   14] = 1'b0;  wr_cycle[   14] = 1'b1;  addr_rom[   14]='h00000038;  wr_data_rom[   14]='h00000062;
    rd_cycle[   15] = 1'b0;  wr_cycle[   15] = 1'b1;  addr_rom[   15]='h0000003c;  wr_data_rom[   15]='h00000159;
    rd_cycle[   16] = 1'b0;  wr_cycle[   16] = 1'b1;  addr_rom[   16]='h00000040;  wr_data_rom[   16]='h00000066;
    rd_cycle[   17] = 1'b0;  wr_cycle[   17] = 1'b1;  addr_rom[   17]='h00000044;  wr_data_rom[   17]='h0000009d;
    rd_cycle[   18] = 1'b0;  wr_cycle[   18] = 1'b1;  addr_rom[   18]='h00000048;  wr_data_rom[   18]='h0000011f;
    rd_cycle[   19] = 1'b0;  wr_cycle[   19] = 1'b1;  addr_rom[   19]='h0000004c;  wr_data_rom[   19]='h00000009;
    rd_cycle[   20] = 1'b0;  wr_cycle[   20] = 1'b1;  addr_rom[   20]='h00000050;  wr_data_rom[   20]='h00000030;
    rd_cycle[   21] = 1'b0;  wr_cycle[   21] = 1'b1;  addr_rom[   21]='h00000054;  wr_data_rom[   21]='h0000007c;
    rd_cycle[   22] = 1'b0;  wr_cycle[   22] = 1'b1;  addr_rom[   22]='h00000058;  wr_data_rom[   22]='h00000006;
    rd_cycle[   23] = 1'b0;  wr_cycle[   23] = 1'b1;  addr_rom[   23]='h0000005c;  wr_data_rom[   23]='h000000fe;
    rd_cycle[   24] = 1'b0;  wr_cycle[   24] = 1'b1;  addr_rom[   24]='h00000060;  wr_data_rom[   24]='h000000e7;
    rd_cycle[   25] = 1'b0;  wr_cycle[   25] = 1'b1;  addr_rom[   25]='h00000064;  wr_data_rom[   25]='h00000026;
    rd_cycle[   26] = 1'b0;  wr_cycle[   26] = 1'b1;  addr_rom[   26]='h00000068;  wr_data_rom[   26]='h0000008d;
    rd_cycle[   27] = 1'b0;  wr_cycle[   27] = 1'b1;  addr_rom[   27]='h0000006c;  wr_data_rom[   27]='h00000072;
    rd_cycle[   28] = 1'b0;  wr_cycle[   28] = 1'b1;  addr_rom[   28]='h00000070;  wr_data_rom[   28]='h000000d4;
    rd_cycle[   29] = 1'b0;  wr_cycle[   29] = 1'b1;  addr_rom[   29]='h00000074;  wr_data_rom[   29]='h0000016e;
    rd_cycle[   30] = 1'b0;  wr_cycle[   30] = 1'b1;  addr_rom[   30]='h00000078;  wr_data_rom[   30]='h00000021;
    rd_cycle[   31] = 1'b0;  wr_cycle[   31] = 1'b1;  addr_rom[   31]='h0000007c;  wr_data_rom[   31]='h00000127;
    rd_cycle[   32] = 1'b0;  wr_cycle[   32] = 1'b1;  addr_rom[   32]='h00000080;  wr_data_rom[   32]='h000000f5;
    rd_cycle[   33] = 1'b0;  wr_cycle[   33] = 1'b1;  addr_rom[   33]='h00000084;  wr_data_rom[   33]='h000000c0;
    rd_cycle[   34] = 1'b0;  wr_cycle[   34] = 1'b1;  addr_rom[   34]='h00000088;  wr_data_rom[   34]='h0000001c;
    rd_cycle[   35] = 1'b0;  wr_cycle[   35] = 1'b1;  addr_rom[   35]='h0000008c;  wr_data_rom[   35]='h00000027;
    rd_cycle[   36] = 1'b0;  wr_cycle[   36] = 1'b1;  addr_rom[   36]='h00000090;  wr_data_rom[   36]='h00000170;
    rd_cycle[   37] = 1'b0;  wr_cycle[   37] = 1'b1;  addr_rom[   37]='h00000094;  wr_data_rom[   37]='h0000015e;
    rd_cycle[   38] = 1'b0;  wr_cycle[   38] = 1'b1;  addr_rom[   38]='h00000098;  wr_data_rom[   38]='h00000036;
    rd_cycle[   39] = 1'b0;  wr_cycle[   39] = 1'b1;  addr_rom[   39]='h0000009c;  wr_data_rom[   39]='h00000098;
    rd_cycle[   40] = 1'b0;  wr_cycle[   40] = 1'b1;  addr_rom[   40]='h000000a0;  wr_data_rom[   40]='h0000005f;
    rd_cycle[   41] = 1'b0;  wr_cycle[   41] = 1'b1;  addr_rom[   41]='h000000a4;  wr_data_rom[   41]='h000000ac;
    rd_cycle[   42] = 1'b0;  wr_cycle[   42] = 1'b1;  addr_rom[   42]='h000000a8;  wr_data_rom[   42]='h00000106;
    rd_cycle[   43] = 1'b0;  wr_cycle[   43] = 1'b1;  addr_rom[   43]='h000000ac;  wr_data_rom[   43]='h0000014b;
    rd_cycle[   44] = 1'b0;  wr_cycle[   44] = 1'b1;  addr_rom[   44]='h000000b0;  wr_data_rom[   44]='h0000001d;
    rd_cycle[   45] = 1'b0;  wr_cycle[   45] = 1'b1;  addr_rom[   45]='h000000b4;  wr_data_rom[   45]='h000000ff;
    rd_cycle[   46] = 1'b0;  wr_cycle[   46] = 1'b1;  addr_rom[   46]='h000000b8;  wr_data_rom[   46]='h000000ec;
    rd_cycle[   47] = 1'b0;  wr_cycle[   47] = 1'b1;  addr_rom[   47]='h000000bc;  wr_data_rom[   47]='h0000001a;
    rd_cycle[   48] = 1'b0;  wr_cycle[   48] = 1'b1;  addr_rom[   48]='h000000c0;  wr_data_rom[   48]='h00000179;
    rd_cycle[   49] = 1'b0;  wr_cycle[   49] = 1'b1;  addr_rom[   49]='h000000c4;  wr_data_rom[   49]='h0000004b;
    rd_cycle[   50] = 1'b0;  wr_cycle[   50] = 1'b1;  addr_rom[   50]='h000000c8;  wr_data_rom[   50]='h000000bf;
    rd_cycle[   51] = 1'b0;  wr_cycle[   51] = 1'b1;  addr_rom[   51]='h000000cc;  wr_data_rom[   51]='h00000017;
    rd_cycle[   52] = 1'b0;  wr_cycle[   52] = 1'b1;  addr_rom[   52]='h000000d0;  wr_data_rom[   52]='h0000018b;
    rd_cycle[   53] = 1'b0;  wr_cycle[   53] = 1'b1;  addr_rom[   53]='h000000d4;  wr_data_rom[   53]='h00000073;
    rd_cycle[   54] = 1'b0;  wr_cycle[   54] = 1'b1;  addr_rom[   54]='h000000d8;  wr_data_rom[   54]='h00000040;
    rd_cycle[   55] = 1'b0;  wr_cycle[   55] = 1'b1;  addr_rom[   55]='h000000dc;  wr_data_rom[   55]='h00000186;
    rd_cycle[   56] = 1'b0;  wr_cycle[   56] = 1'b1;  addr_rom[   56]='h000000e0;  wr_data_rom[   56]='h00000029;
    rd_cycle[   57] = 1'b0;  wr_cycle[   57] = 1'b1;  addr_rom[   57]='h000000e4;  wr_data_rom[   57]='h0000013e;
    rd_cycle[   58] = 1'b0;  wr_cycle[   58] = 1'b1;  addr_rom[   58]='h000000e8;  wr_data_rom[   58]='h000000d9;
    rd_cycle[   59] = 1'b0;  wr_cycle[   59] = 1'b1;  addr_rom[   59]='h000000ec;  wr_data_rom[   59]='h00000046;
    rd_cycle[   60] = 1'b0;  wr_cycle[   60] = 1'b1;  addr_rom[   60]='h000000f0;  wr_data_rom[   60]='h000000c1;
    rd_cycle[   61] = 1'b0;  wr_cycle[   61] = 1'b1;  addr_rom[   61]='h000000f4;  wr_data_rom[   61]='h000000ad;
    rd_cycle[   62] = 1'b0;  wr_cycle[   62] = 1'b1;  addr_rom[   62]='h000000f8;  wr_data_rom[   62]='h00000178;
    rd_cycle[   63] = 1'b0;  wr_cycle[   63] = 1'b1;  addr_rom[   63]='h000000fc;  wr_data_rom[   63]='h000000fc;
    rd_cycle[   64] = 1'b0;  wr_cycle[   64] = 1'b1;  addr_rom[   64]='h00000100;  wr_data_rom[   64]='h0000015e;
    rd_cycle[   65] = 1'b0;  wr_cycle[   65] = 1'b1;  addr_rom[   65]='h00000104;  wr_data_rom[   65]='h00000011;
    rd_cycle[   66] = 1'b0;  wr_cycle[   66] = 1'b1;  addr_rom[   66]='h00000108;  wr_data_rom[   66]='h00000090;
    rd_cycle[   67] = 1'b0;  wr_cycle[   67] = 1'b1;  addr_rom[   67]='h0000010c;  wr_data_rom[   67]='h0000011e;
    rd_cycle[   68] = 1'b0;  wr_cycle[   68] = 1'b1;  addr_rom[   68]='h00000110;  wr_data_rom[   68]='h000000c8;
    rd_cycle[   69] = 1'b0;  wr_cycle[   69] = 1'b1;  addr_rom[   69]='h00000114;  wr_data_rom[   69]='h0000007d;
    rd_cycle[   70] = 1'b0;  wr_cycle[   70] = 1'b1;  addr_rom[   70]='h00000118;  wr_data_rom[   70]='h0000002a;
    rd_cycle[   71] = 1'b0;  wr_cycle[   71] = 1'b1;  addr_rom[   71]='h0000011c;  wr_data_rom[   71]='h0000008b;
    rd_cycle[   72] = 1'b0;  wr_cycle[   72] = 1'b1;  addr_rom[   72]='h00000120;  wr_data_rom[   72]='h0000008f;
    rd_cycle[   73] = 1'b0;  wr_cycle[   73] = 1'b1;  addr_rom[   73]='h00000124;  wr_data_rom[   73]='h000000b5;
    rd_cycle[   74] = 1'b0;  wr_cycle[   74] = 1'b1;  addr_rom[   74]='h00000128;  wr_data_rom[   74]='h00000026;
    rd_cycle[   75] = 1'b0;  wr_cycle[   75] = 1'b1;  addr_rom[   75]='h0000012c;  wr_data_rom[   75]='h00000163;
    rd_cycle[   76] = 1'b0;  wr_cycle[   76] = 1'b1;  addr_rom[   76]='h00000130;  wr_data_rom[   76]='h00000156;
    rd_cycle[   77] = 1'b0;  wr_cycle[   77] = 1'b1;  addr_rom[   77]='h00000134;  wr_data_rom[   77]='h000000cb;
    rd_cycle[   78] = 1'b0;  wr_cycle[   78] = 1'b1;  addr_rom[   78]='h00000138;  wr_data_rom[   78]='h00000173;
    rd_cycle[   79] = 1'b0;  wr_cycle[   79] = 1'b1;  addr_rom[   79]='h0000013c;  wr_data_rom[   79]='h000000c0;
    rd_cycle[   80] = 1'b0;  wr_cycle[   80] = 1'b1;  addr_rom[   80]='h00000140;  wr_data_rom[   80]='h0000018d;
    rd_cycle[   81] = 1'b0;  wr_cycle[   81] = 1'b1;  addr_rom[   81]='h00000144;  wr_data_rom[   81]='h00000113;
    rd_cycle[   82] = 1'b0;  wr_cycle[   82] = 1'b1;  addr_rom[   82]='h00000148;  wr_data_rom[   82]='h000000d7;
    rd_cycle[   83] = 1'b0;  wr_cycle[   83] = 1'b1;  addr_rom[   83]='h0000014c;  wr_data_rom[   83]='h00000153;
    rd_cycle[   84] = 1'b0;  wr_cycle[   84] = 1'b1;  addr_rom[   84]='h00000150;  wr_data_rom[   84]='h00000070;
    rd_cycle[   85] = 1'b0;  wr_cycle[   85] = 1'b1;  addr_rom[   85]='h00000154;  wr_data_rom[   85]='h0000016d;
    rd_cycle[   86] = 1'b0;  wr_cycle[   86] = 1'b1;  addr_rom[   86]='h00000158;  wr_data_rom[   86]='h00000022;
    rd_cycle[   87] = 1'b0;  wr_cycle[   87] = 1'b1;  addr_rom[   87]='h0000015c;  wr_data_rom[   87]='h00000029;
    rd_cycle[   88] = 1'b0;  wr_cycle[   88] = 1'b1;  addr_rom[   88]='h00000160;  wr_data_rom[   88]='h000000f7;
    rd_cycle[   89] = 1'b0;  wr_cycle[   89] = 1'b1;  addr_rom[   89]='h00000164;  wr_data_rom[   89]='h00000057;
    rd_cycle[   90] = 1'b0;  wr_cycle[   90] = 1'b1;  addr_rom[   90]='h00000168;  wr_data_rom[   90]='h000000b0;
    rd_cycle[   91] = 1'b0;  wr_cycle[   91] = 1'b1;  addr_rom[   91]='h0000016c;  wr_data_rom[   91]='h000000c3;
    rd_cycle[   92] = 1'b0;  wr_cycle[   92] = 1'b1;  addr_rom[   92]='h00000170;  wr_data_rom[   92]='h0000014d;
    rd_cycle[   93] = 1'b0;  wr_cycle[   93] = 1'b1;  addr_rom[   93]='h00000174;  wr_data_rom[   93]='h0000001b;
    rd_cycle[   94] = 1'b0;  wr_cycle[   94] = 1'b1;  addr_rom[   94]='h00000178;  wr_data_rom[   94]='h0000015a;
    rd_cycle[   95] = 1'b0;  wr_cycle[   95] = 1'b1;  addr_rom[   95]='h0000017c;  wr_data_rom[   95]='h0000002b;
    rd_cycle[   96] = 1'b0;  wr_cycle[   96] = 1'b1;  addr_rom[   96]='h00000180;  wr_data_rom[   96]='h00000177;
    rd_cycle[   97] = 1'b0;  wr_cycle[   97] = 1'b1;  addr_rom[   97]='h00000184;  wr_data_rom[   97]='h00000138;
    rd_cycle[   98] = 1'b0;  wr_cycle[   98] = 1'b1;  addr_rom[   98]='h00000188;  wr_data_rom[   98]='h00000116;
    rd_cycle[   99] = 1'b0;  wr_cycle[   99] = 1'b1;  addr_rom[   99]='h0000018c;  wr_data_rom[   99]='h00000173;
    // 300 random read and write cycles
    rd_cycle[  100] = 1'b0;  wr_cycle[  100] = 1'b1;  addr_rom[  100]='h000000f8;  wr_data_rom[  100]='h0000011b;
    rd_cycle[  101] = 1'b1;  wr_cycle[  101] = 1'b0;  addr_rom[  101]='h00000120;  wr_data_rom[  101]='h00000000;
    rd_cycle[  102] = 1'b0;  wr_cycle[  102] = 1'b1;  addr_rom[  102]='h000000e4;  wr_data_rom[  102]='h00000084;
    rd_cycle[  103] = 1'b0;  wr_cycle[  103] = 1'b1;  addr_rom[  103]='h00000178;  wr_data_rom[  103]='h00000085;
    rd_cycle[  104] = 1'b0;  wr_cycle[  104] = 1'b1;  addr_rom[  104]='h000000d0;  wr_data_rom[  104]='h000000b0;
    rd_cycle[  105] = 1'b1;  wr_cycle[  105] = 1'b0;  addr_rom[  105]='h00000168;  wr_data_rom[  105]='h00000000;
    rd_cycle[  106] = 1'b1;  wr_cycle[  106] = 1'b0;  addr_rom[  106]='h00000070;  wr_data_rom[  106]='h00000000;
    rd_cycle[  107] = 1'b0;  wr_cycle[  107] = 1'b1;  addr_rom[  107]='h0000014c;  wr_data_rom[  107]='h00000056;
    rd_cycle[  108] = 1'b1;  wr_cycle[  108] = 1'b0;  addr_rom[  108]='h00000050;  wr_data_rom[  108]='h00000000;
    rd_cycle[  109] = 1'b1;  wr_cycle[  109] = 1'b0;  addr_rom[  109]='h00000168;  wr_data_rom[  109]='h00000000;
    rd_cycle[  110] = 1'b1;  wr_cycle[  110] = 1'b0;  addr_rom[  110]='h0000018c;  wr_data_rom[  110]='h00000000;
    rd_cycle[  111] = 1'b0;  wr_cycle[  111] = 1'b1;  addr_rom[  111]='h00000120;  wr_data_rom[  111]='h0000009e;
    rd_cycle[  112] = 1'b1;  wr_cycle[  112] = 1'b0;  addr_rom[  112]='h0000011c;  wr_data_rom[  112]='h00000000;
    rd_cycle[  113] = 1'b1;  wr_cycle[  113] = 1'b0;  addr_rom[  113]='h00000024;  wr_data_rom[  113]='h00000000;
    rd_cycle[  114] = 1'b1;  wr_cycle[  114] = 1'b0;  addr_rom[  114]='h000000a4;  wr_data_rom[  114]='h00000000;
    rd_cycle[  115] = 1'b1;  wr_cycle[  115] = 1'b0;  addr_rom[  115]='h00000098;  wr_data_rom[  115]='h00000000;
    rd_cycle[  116] = 1'b0;  wr_cycle[  116] = 1'b1;  addr_rom[  116]='h00000108;  wr_data_rom[  116]='h00000033;
    rd_cycle[  117] = 1'b1;  wr_cycle[  117] = 1'b0;  addr_rom[  117]='h00000094;  wr_data_rom[  117]='h00000000;
    rd_cycle[  118] = 1'b1;  wr_cycle[  118] = 1'b0;  addr_rom[  118]='h00000160;  wr_data_rom[  118]='h00000000;
    rd_cycle[  119] = 1'b1;  wr_cycle[  119] = 1'b0;  addr_rom[  119]='h00000088;  wr_data_rom[  119]='h00000000;
    rd_cycle[  120] = 1'b0;  wr_cycle[  120] = 1'b1;  addr_rom[  120]='h00000110;  wr_data_rom[  120]='h00000172;
    rd_cycle[  121] = 1'b0;  wr_cycle[  121] = 1'b1;  addr_rom[  121]='h00000080;  wr_data_rom[  121]='h0000016e;
    rd_cycle[  122] = 1'b1;  wr_cycle[  122] = 1'b0;  addr_rom[  122]='h00000180;  wr_data_rom[  122]='h00000000;
    rd_cycle[  123] = 1'b0;  wr_cycle[  123] = 1'b1;  addr_rom[  123]='h00000150;  wr_data_rom[  123]='h00000090;
    rd_cycle[  124] = 1'b1;  wr_cycle[  124] = 1'b0;  addr_rom[  124]='h000000b8;  wr_data_rom[  124]='h00000000;
    rd_cycle[  125] = 1'b0;  wr_cycle[  125] = 1'b1;  addr_rom[  125]='h000000d8;  wr_data_rom[  125]='h00000011;
    rd_cycle[  126] = 1'b1;  wr_cycle[  126] = 1'b0;  addr_rom[  126]='h0000012c;  wr_data_rom[  126]='h00000000;
    rd_cycle[  127] = 1'b0;  wr_cycle[  127] = 1'b1;  addr_rom[  127]='h00000068;  wr_data_rom[  127]='h0000005d;
    rd_cycle[  128] = 1'b1;  wr_cycle[  128] = 1'b0;  addr_rom[  128]='h00000140;  wr_data_rom[  128]='h00000000;
    rd_cycle[  129] = 1'b1;  wr_cycle[  129] = 1'b0;  addr_rom[  129]='h00000158;  wr_data_rom[  129]='h00000000;
    rd_cycle[  130] = 1'b1;  wr_cycle[  130] = 1'b0;  addr_rom[  130]='h00000048;  wr_data_rom[  130]='h00000000;
    rd_cycle[  131] = 1'b0;  wr_cycle[  131] = 1'b1;  addr_rom[  131]='h00000140;  wr_data_rom[  131]='h0000007a;
    rd_cycle[  132] = 1'b1;  wr_cycle[  132] = 1'b0;  addr_rom[  132]='h00000030;  wr_data_rom[  132]='h00000000;
    rd_cycle[  133] = 1'b1;  wr_cycle[  133] = 1'b0;  addr_rom[  133]='h00000074;  wr_data_rom[  133]='h00000000;
    rd_cycle[  134] = 1'b0;  wr_cycle[  134] = 1'b1;  addr_rom[  134]='h000000f4;  wr_data_rom[  134]='h0000013f;
    rd_cycle[  135] = 1'b1;  wr_cycle[  135] = 1'b0;  addr_rom[  135]='h00000048;  wr_data_rom[  135]='h00000000;
    rd_cycle[  136] = 1'b0;  wr_cycle[  136] = 1'b1;  addr_rom[  136]='h000000a4;  wr_data_rom[  136]='h0000015d;
    rd_cycle[  137] = 1'b1;  wr_cycle[  137] = 1'b0;  addr_rom[  137]='h00000130;  wr_data_rom[  137]='h00000000;
    rd_cycle[  138] = 1'b1;  wr_cycle[  138] = 1'b0;  addr_rom[  138]='h000000c0;  wr_data_rom[  138]='h00000000;
    rd_cycle[  139] = 1'b1;  wr_cycle[  139] = 1'b0;  addr_rom[  139]='h000000e4;  wr_data_rom[  139]='h00000000;
    rd_cycle[  140] = 1'b1;  wr_cycle[  140] = 1'b0;  addr_rom[  140]='h0000013c;  wr_data_rom[  140]='h00000000;
    rd_cycle[  141] = 1'b1;  wr_cycle[  141] = 1'b0;  addr_rom[  141]='h00000114;  wr_data_rom[  141]='h00000000;
    rd_cycle[  142] = 1'b1;  wr_cycle[  142] = 1'b0;  addr_rom[  142]='h000000f0;  wr_data_rom[  142]='h00000000;
    rd_cycle[  143] = 1'b0;  wr_cycle[  143] = 1'b1;  addr_rom[  143]='h00000140;  wr_data_rom[  143]='h00000009;
    rd_cycle[  144] = 1'b0;  wr_cycle[  144] = 1'b1;  addr_rom[  144]='h0000010c;  wr_data_rom[  144]='h00000180;
    rd_cycle[  145] = 1'b1;  wr_cycle[  145] = 1'b0;  addr_rom[  145]='h0000013c;  wr_data_rom[  145]='h00000000;
    rd_cycle[  146] = 1'b0;  wr_cycle[  146] = 1'b1;  addr_rom[  146]='h000000b8;  wr_data_rom[  146]='h0000004c;
    rd_cycle[  147] = 1'b0;  wr_cycle[  147] = 1'b1;  addr_rom[  147]='h00000048;  wr_data_rom[  147]='h00000065;
    rd_cycle[  148] = 1'b1;  wr_cycle[  148] = 1'b0;  addr_rom[  148]='h000000e0;  wr_data_rom[  148]='h00000000;
    rd_cycle[  149] = 1'b1;  wr_cycle[  149] = 1'b0;  addr_rom[  149]='h0000005c;  wr_data_rom[  149]='h00000000;
    rd_cycle[  150] = 1'b0;  wr_cycle[  150] = 1'b1;  addr_rom[  150]='h00000064;  wr_data_rom[  150]='h000000a1;
    rd_cycle[  151] = 1'b1;  wr_cycle[  151] = 1'b0;  addr_rom[  151]='h00000064;  wr_data_rom[  151]='h00000000;
    rd_cycle[  152] = 1'b1;  wr_cycle[  152] = 1'b0;  addr_rom[  152]='h0000015c;  wr_data_rom[  152]='h00000000;
    rd_cycle[  153] = 1'b0;  wr_cycle[  153] = 1'b1;  addr_rom[  153]='h000000a8;  wr_data_rom[  153]='h00000045;
    rd_cycle[  154] = 1'b0;  wr_cycle[  154] = 1'b1;  addr_rom[  154]='h00000020;  wr_data_rom[  154]='h00000085;
    rd_cycle[  155] = 1'b1;  wr_cycle[  155] = 1'b0;  addr_rom[  155]='h00000050;  wr_data_rom[  155]='h00000000;
    rd_cycle[  156] = 1'b1;  wr_cycle[  156] = 1'b0;  addr_rom[  156]='h000000a0;  wr_data_rom[  156]='h00000000;
    rd_cycle[  157] = 1'b1;  wr_cycle[  157] = 1'b0;  addr_rom[  157]='h000000bc;  wr_data_rom[  157]='h00000000;
    rd_cycle[  158] = 1'b1;  wr_cycle[  158] = 1'b0;  addr_rom[  158]='h00000130;  wr_data_rom[  158]='h00000000;
    rd_cycle[  159] = 1'b1;  wr_cycle[  159] = 1'b0;  addr_rom[  159]='h000000f4;  wr_data_rom[  159]='h00000000;
    rd_cycle[  160] = 1'b1;  wr_cycle[  160] = 1'b0;  addr_rom[  160]='h00000020;  wr_data_rom[  160]='h00000000;
    rd_cycle[  161] = 1'b0;  wr_cycle[  161] = 1'b1;  addr_rom[  161]='h000000ac;  wr_data_rom[  161]='h0000007f;
    rd_cycle[  162] = 1'b1;  wr_cycle[  162] = 1'b0;  addr_rom[  162]='h0000018c;  wr_data_rom[  162]='h00000000;
    rd_cycle[  163] = 1'b1;  wr_cycle[  163] = 1'b0;  addr_rom[  163]='h00000020;  wr_data_rom[  163]='h00000000;
    rd_cycle[  164] = 1'b0;  wr_cycle[  164] = 1'b1;  addr_rom[  164]='h00000110;  wr_data_rom[  164]='h0000016d;
    rd_cycle[  165] = 1'b1;  wr_cycle[  165] = 1'b0;  addr_rom[  165]='h00000068;  wr_data_rom[  165]='h00000000;
    rd_cycle[  166] = 1'b0;  wr_cycle[  166] = 1'b1;  addr_rom[  166]='h000000dc;  wr_data_rom[  166]='h00000077;
    rd_cycle[  167] = 1'b1;  wr_cycle[  167] = 1'b0;  addr_rom[  167]='h00000104;  wr_data_rom[  167]='h00000000;
    rd_cycle[  168] = 1'b1;  wr_cycle[  168] = 1'b0;  addr_rom[  168]='h00000140;  wr_data_rom[  168]='h00000000;
    rd_cycle[  169] = 1'b0;  wr_cycle[  169] = 1'b1;  addr_rom[  169]='h00000094;  wr_data_rom[  169]='h0000011e;
    rd_cycle[  170] = 1'b0;  wr_cycle[  170] = 1'b1;  addr_rom[  170]='h00000024;  wr_data_rom[  170]='h00000068;
    rd_cycle[  171] = 1'b1;  wr_cycle[  171] = 1'b0;  addr_rom[  171]='h00000108;  wr_data_rom[  171]='h00000000;
    rd_cycle[  172] = 1'b0;  wr_cycle[  172] = 1'b1;  addr_rom[  172]='h000000f8;  wr_data_rom[  172]='h00000062;
    rd_cycle[  173] = 1'b1;  wr_cycle[  173] = 1'b0;  addr_rom[  173]='h00000174;  wr_data_rom[  173]='h00000000;
    rd_cycle[  174] = 1'b0;  wr_cycle[  174] = 1'b1;  addr_rom[  174]='h0000016c;  wr_data_rom[  174]='h0000000e;
    rd_cycle[  175] = 1'b1;  wr_cycle[  175] = 1'b0;  addr_rom[  175]='h00000178;  wr_data_rom[  175]='h00000000;
    rd_cycle[  176] = 1'b1;  wr_cycle[  176] = 1'b0;  addr_rom[  176]='h00000024;  wr_data_rom[  176]='h00000000;
    rd_cycle[  177] = 1'b1;  wr_cycle[  177] = 1'b0;  addr_rom[  177]='h00000104;  wr_data_rom[  177]='h00000000;
    rd_cycle[  178] = 1'b0;  wr_cycle[  178] = 1'b1;  addr_rom[  178]='h00000084;  wr_data_rom[  178]='h00000063;
    rd_cycle[  179] = 1'b1;  wr_cycle[  179] = 1'b0;  addr_rom[  179]='h000000ac;  wr_data_rom[  179]='h00000000;
    rd_cycle[  180] = 1'b1;  wr_cycle[  180] = 1'b0;  addr_rom[  180]='h00000080;  wr_data_rom[  180]='h00000000;
    rd_cycle[  181] = 1'b1;  wr_cycle[  181] = 1'b0;  addr_rom[  181]='h0000008c;  wr_data_rom[  181]='h00000000;
    rd_cycle[  182] = 1'b1;  wr_cycle[  182] = 1'b0;  addr_rom[  182]='h000000e4;  wr_data_rom[  182]='h00000000;
    rd_cycle[  183] = 1'b0;  wr_cycle[  183] = 1'b1;  addr_rom[  183]='h00000060;  wr_data_rom[  183]='h00000094;
    rd_cycle[  184] = 1'b0;  wr_cycle[  184] = 1'b1;  addr_rom[  184]='h000000ac;  wr_data_rom[  184]='h000000e8;
    rd_cycle[  185] = 1'b1;  wr_cycle[  185] = 1'b0;  addr_rom[  185]='h000000ec;  wr_data_rom[  185]='h00000000;
    rd_cycle[  186] = 1'b0;  wr_cycle[  186] = 1'b1;  addr_rom[  186]='h00000058;  wr_data_rom[  186]='h00000010;
    rd_cycle[  187] = 1'b1;  wr_cycle[  187] = 1'b0;  addr_rom[  187]='h00000050;  wr_data_rom[  187]='h00000000;
    rd_cycle[  188] = 1'b1;  wr_cycle[  188] = 1'b0;  addr_rom[  188]='h00000078;  wr_data_rom[  188]='h00000000;
    rd_cycle[  189] = 1'b0;  wr_cycle[  189] = 1'b1;  addr_rom[  189]='h000000fc;  wr_data_rom[  189]='h0000012b;
    rd_cycle[  190] = 1'b0;  wr_cycle[  190] = 1'b1;  addr_rom[  190]='h000000e0;  wr_data_rom[  190]='h00000065;
    rd_cycle[  191] = 1'b1;  wr_cycle[  191] = 1'b0;  addr_rom[  191]='h00000168;  wr_data_rom[  191]='h00000000;
    rd_cycle[  192] = 1'b1;  wr_cycle[  192] = 1'b0;  addr_rom[  192]='h00000148;  wr_data_rom[  192]='h00000000;
    rd_cycle[  193] = 1'b0;  wr_cycle[  193] = 1'b1;  addr_rom[  193]='h00000168;  wr_data_rom[  193]='h00000091;
    rd_cycle[  194] = 1'b0;  wr_cycle[  194] = 1'b1;  addr_rom[  194]='h00000070;  wr_data_rom[  194]='h0000013f;
    rd_cycle[  195] = 1'b0;  wr_cycle[  195] = 1'b1;  addr_rom[  195]='h00000050;  wr_data_rom[  195]='h00000113;
    rd_cycle[  196] = 1'b1;  wr_cycle[  196] = 1'b0;  addr_rom[  196]='h00000060;  wr_data_rom[  196]='h00000000;
    rd_cycle[  197] = 1'b0;  wr_cycle[  197] = 1'b1;  addr_rom[  197]='h000000e0;  wr_data_rom[  197]='h000000f9;
    rd_cycle[  198] = 1'b0;  wr_cycle[  198] = 1'b1;  addr_rom[  198]='h000000bc;  wr_data_rom[  198]='h00000173;
    rd_cycle[  199] = 1'b1;  wr_cycle[  199] = 1'b0;  addr_rom[  199]='h00000068;  wr_data_rom[  199]='h00000000;
    rd_cycle[  200] = 1'b1;  wr_cycle[  200] = 1'b0;  addr_rom[  200]='h00000014;  wr_data_rom[  200]='h00000000;
    rd_cycle[  201] = 1'b1;  wr_cycle[  201] = 1'b0;  addr_rom[  201]='h00000018;  wr_data_rom[  201]='h00000000;
    rd_cycle[  202] = 1'b1;  wr_cycle[  202] = 1'b0;  addr_rom[  202]='h000000cc;  wr_data_rom[  202]='h00000000;
    rd_cycle[  203] = 1'b0;  wr_cycle[  203] = 1'b1;  addr_rom[  203]='h000000f8;  wr_data_rom[  203]='h00000047;
    rd_cycle[  204] = 1'b1;  wr_cycle[  204] = 1'b0;  addr_rom[  204]='h00000154;  wr_data_rom[  204]='h00000000;
    rd_cycle[  205] = 1'b1;  wr_cycle[  205] = 1'b0;  addr_rom[  205]='h00000008;  wr_data_rom[  205]='h00000000;
    rd_cycle[  206] = 1'b0;  wr_cycle[  206] = 1'b1;  addr_rom[  206]='h00000030;  wr_data_rom[  206]='h00000147;
    rd_cycle[  207] = 1'b1;  wr_cycle[  207] = 1'b0;  addr_rom[  207]='h00000058;  wr_data_rom[  207]='h00000000;
    rd_cycle[  208] = 1'b1;  wr_cycle[  208] = 1'b0;  addr_rom[  208]='h00000040;  wr_data_rom[  208]='h00000000;
    rd_cycle[  209] = 1'b0;  wr_cycle[  209] = 1'b1;  addr_rom[  209]='h00000180;  wr_data_rom[  209]='h000000c1;
    rd_cycle[  210] = 1'b1;  wr_cycle[  210] = 1'b0;  addr_rom[  210]='h00000074;  wr_data_rom[  210]='h00000000;
    rd_cycle[  211] = 1'b0;  wr_cycle[  211] = 1'b1;  addr_rom[  211]='h00000120;  wr_data_rom[  211]='h00000183;
    rd_cycle[  212] = 1'b0;  wr_cycle[  212] = 1'b1;  addr_rom[  212]='h00000050;  wr_data_rom[  212]='h000000f0;
    rd_cycle[  213] = 1'b1;  wr_cycle[  213] = 1'b0;  addr_rom[  213]='h00000020;  wr_data_rom[  213]='h00000000;
    rd_cycle[  214] = 1'b0;  wr_cycle[  214] = 1'b1;  addr_rom[  214]='h00000140;  wr_data_rom[  214]='h00000142;
    rd_cycle[  215] = 1'b1;  wr_cycle[  215] = 1'b0;  addr_rom[  215]='h00000080;  wr_data_rom[  215]='h00000000;
    rd_cycle[  216] = 1'b0;  wr_cycle[  216] = 1'b1;  addr_rom[  216]='h000000a8;  wr_data_rom[  216]='h00000060;
    rd_cycle[  217] = 1'b0;  wr_cycle[  217] = 1'b1;  addr_rom[  217]='h000000c0;  wr_data_rom[  217]='h00000178;
    rd_cycle[  218] = 1'b1;  wr_cycle[  218] = 1'b0;  addr_rom[  218]='h000000c4;  wr_data_rom[  218]='h00000000;
    rd_cycle[  219] = 1'b0;  wr_cycle[  219] = 1'b1;  addr_rom[  219]='h00000114;  wr_data_rom[  219]='h000000ce;
    rd_cycle[  220] = 1'b1;  wr_cycle[  220] = 1'b0;  addr_rom[  220]='h0000005c;  wr_data_rom[  220]='h00000000;
    rd_cycle[  221] = 1'b0;  wr_cycle[  221] = 1'b1;  addr_rom[  221]='h000000ac;  wr_data_rom[  221]='h0000014d;
    rd_cycle[  222] = 1'b1;  wr_cycle[  222] = 1'b0;  addr_rom[  222]='h000000dc;  wr_data_rom[  222]='h00000000;
    rd_cycle[  223] = 1'b0;  wr_cycle[  223] = 1'b1;  addr_rom[  223]='h00000038;  wr_data_rom[  223]='h00000015;
    rd_cycle[  224] = 1'b1;  wr_cycle[  224] = 1'b0;  addr_rom[  224]='h000000a4;  wr_data_rom[  224]='h00000000;
    rd_cycle[  225] = 1'b0;  wr_cycle[  225] = 1'b1;  addr_rom[  225]='h00000144;  wr_data_rom[  225]='h000000a1;
    rd_cycle[  226] = 1'b0;  wr_cycle[  226] = 1'b1;  addr_rom[  226]='h00000050;  wr_data_rom[  226]='h0000011c;
    rd_cycle[  227] = 1'b0;  wr_cycle[  227] = 1'b1;  addr_rom[  227]='h00000150;  wr_data_rom[  227]='h000000f9;
    rd_cycle[  228] = 1'b0;  wr_cycle[  228] = 1'b1;  addr_rom[  228]='h00000154;  wr_data_rom[  228]='h0000014d;
    rd_cycle[  229] = 1'b1;  wr_cycle[  229] = 1'b0;  addr_rom[  229]='h000000c4;  wr_data_rom[  229]='h00000000;
    rd_cycle[  230] = 1'b0;  wr_cycle[  230] = 1'b1;  addr_rom[  230]='h0000002c;  wr_data_rom[  230]='h00000186;
    rd_cycle[  231] = 1'b1;  wr_cycle[  231] = 1'b0;  addr_rom[  231]='h00000104;  wr_data_rom[  231]='h00000000;
    rd_cycle[  232] = 1'b0;  wr_cycle[  232] = 1'b1;  addr_rom[  232]='h00000110;  wr_data_rom[  232]='h0000015e;
    rd_cycle[  233] = 1'b0;  wr_cycle[  233] = 1'b1;  addr_rom[  233]='h00000028;  wr_data_rom[  233]='h000000a5;
    rd_cycle[  234] = 1'b0;  wr_cycle[  234] = 1'b1;  addr_rom[  234]='h00000028;  wr_data_rom[  234]='h00000148;
    rd_cycle[  235] = 1'b1;  wr_cycle[  235] = 1'b0;  addr_rom[  235]='h00000068;  wr_data_rom[  235]='h00000000;
    rd_cycle[  236] = 1'b0;  wr_cycle[  236] = 1'b1;  addr_rom[  236]='h000000c4;  wr_data_rom[  236]='h0000003e;
    rd_cycle[  237] = 1'b1;  wr_cycle[  237] = 1'b0;  addr_rom[  237]='h000000bc;  wr_data_rom[  237]='h00000000;
    rd_cycle[  238] = 1'b0;  wr_cycle[  238] = 1'b1;  addr_rom[  238]='h00000164;  wr_data_rom[  238]='h000000bf;
    rd_cycle[  239] = 1'b1;  wr_cycle[  239] = 1'b0;  addr_rom[  239]='h00000038;  wr_data_rom[  239]='h00000000;
    rd_cycle[  240] = 1'b1;  wr_cycle[  240] = 1'b0;  addr_rom[  240]='h00000078;  wr_data_rom[  240]='h00000000;
    rd_cycle[  241] = 1'b1;  wr_cycle[  241] = 1'b0;  addr_rom[  241]='h00000110;  wr_data_rom[  241]='h00000000;
    rd_cycle[  242] = 1'b0;  wr_cycle[  242] = 1'b1;  addr_rom[  242]='h0000003c;  wr_data_rom[  242]='h00000100;
    rd_cycle[  243] = 1'b0;  wr_cycle[  243] = 1'b1;  addr_rom[  243]='h00000160;  wr_data_rom[  243]='h000000ce;
    rd_cycle[  244] = 1'b0;  wr_cycle[  244] = 1'b1;  addr_rom[  244]='h00000050;  wr_data_rom[  244]='h0000011b;
    rd_cycle[  245] = 1'b0;  wr_cycle[  245] = 1'b1;  addr_rom[  245]='h00000078;  wr_data_rom[  245]='h00000029;
    rd_cycle[  246] = 1'b1;  wr_cycle[  246] = 1'b0;  addr_rom[  246]='h00000078;  wr_data_rom[  246]='h00000000;
    rd_cycle[  247] = 1'b0;  wr_cycle[  247] = 1'b1;  addr_rom[  247]='h00000040;  wr_data_rom[  247]='h00000028;
    rd_cycle[  248] = 1'b0;  wr_cycle[  248] = 1'b1;  addr_rom[  248]='h000000fc;  wr_data_rom[  248]='h00000098;
    rd_cycle[  249] = 1'b0;  wr_cycle[  249] = 1'b1;  addr_rom[  249]='h00000090;  wr_data_rom[  249]='h00000141;
    rd_cycle[  250] = 1'b0;  wr_cycle[  250] = 1'b1;  addr_rom[  250]='h0000001c;  wr_data_rom[  250]='h00000055;
    rd_cycle[  251] = 1'b0;  wr_cycle[  251] = 1'b1;  addr_rom[  251]='h00000070;  wr_data_rom[  251]='h0000002e;
    rd_cycle[  252] = 1'b1;  wr_cycle[  252] = 1'b0;  addr_rom[  252]='h000000e4;  wr_data_rom[  252]='h00000000;
    rd_cycle[  253] = 1'b0;  wr_cycle[  253] = 1'b1;  addr_rom[  253]='h0000012c;  wr_data_rom[  253]='h000000aa;
    rd_cycle[  254] = 1'b1;  wr_cycle[  254] = 1'b0;  addr_rom[  254]='h00000088;  wr_data_rom[  254]='h00000000;
    rd_cycle[  255] = 1'b1;  wr_cycle[  255] = 1'b0;  addr_rom[  255]='h00000030;  wr_data_rom[  255]='h00000000;
    rd_cycle[  256] = 1'b0;  wr_cycle[  256] = 1'b1;  addr_rom[  256]='h00000004;  wr_data_rom[  256]='h0000011d;
    rd_cycle[  257] = 1'b0;  wr_cycle[  257] = 1'b1;  addr_rom[  257]='h00000064;  wr_data_rom[  257]='h00000115;
    rd_cycle[  258] = 1'b0;  wr_cycle[  258] = 1'b1;  addr_rom[  258]='h00000090;  wr_data_rom[  258]='h0000009b;
    rd_cycle[  259] = 1'b0;  wr_cycle[  259] = 1'b1;  addr_rom[  259]='h000000fc;  wr_data_rom[  259]='h0000001d;
    rd_cycle[  260] = 1'b1;  wr_cycle[  260] = 1'b0;  addr_rom[  260]='h0000004c;  wr_data_rom[  260]='h00000000;
    rd_cycle[  261] = 1'b0;  wr_cycle[  261] = 1'b1;  addr_rom[  261]='h00000108;  wr_data_rom[  261]='h00000054;
    rd_cycle[  262] = 1'b1;  wr_cycle[  262] = 1'b0;  addr_rom[  262]='h00000078;  wr_data_rom[  262]='h00000000;
    rd_cycle[  263] = 1'b0;  wr_cycle[  263] = 1'b1;  addr_rom[  263]='h0000013c;  wr_data_rom[  263]='h00000126;
    rd_cycle[  264] = 1'b0;  wr_cycle[  264] = 1'b1;  addr_rom[  264]='h00000118;  wr_data_rom[  264]='h00000173;
    rd_cycle[  265] = 1'b1;  wr_cycle[  265] = 1'b0;  addr_rom[  265]='h00000028;  wr_data_rom[  265]='h00000000;
    rd_cycle[  266] = 1'b1;  wr_cycle[  266] = 1'b0;  addr_rom[  266]='h00000004;  wr_data_rom[  266]='h00000000;
    rd_cycle[  267] = 1'b1;  wr_cycle[  267] = 1'b0;  addr_rom[  267]='h00000080;  wr_data_rom[  267]='h00000000;
    rd_cycle[  268] = 1'b1;  wr_cycle[  268] = 1'b0;  addr_rom[  268]='h00000124;  wr_data_rom[  268]='h00000000;
    rd_cycle[  269] = 1'b0;  wr_cycle[  269] = 1'b1;  addr_rom[  269]='h000000f8;  wr_data_rom[  269]='h000000b6;
    rd_cycle[  270] = 1'b0;  wr_cycle[  270] = 1'b1;  addr_rom[  270]='h00000114;  wr_data_rom[  270]='h000000fa;
    rd_cycle[  271] = 1'b0;  wr_cycle[  271] = 1'b1;  addr_rom[  271]='h000000e4;  wr_data_rom[  271]='h000000ea;
    rd_cycle[  272] = 1'b1;  wr_cycle[  272] = 1'b0;  addr_rom[  272]='h00000094;  wr_data_rom[  272]='h00000000;
    rd_cycle[  273] = 1'b1;  wr_cycle[  273] = 1'b0;  addr_rom[  273]='h00000164;  wr_data_rom[  273]='h00000000;
    rd_cycle[  274] = 1'b0;  wr_cycle[  274] = 1'b1;  addr_rom[  274]='h00000064;  wr_data_rom[  274]='h00000161;
    rd_cycle[  275] = 1'b0;  wr_cycle[  275] = 1'b1;  addr_rom[  275]='h000000b8;  wr_data_rom[  275]='h0000001f;
    rd_cycle[  276] = 1'b0;  wr_cycle[  276] = 1'b1;  addr_rom[  276]='h0000003c;  wr_data_rom[  276]='h000000b2;
    rd_cycle[  277] = 1'b0;  wr_cycle[  277] = 1'b1;  addr_rom[  277]='h000000d8;  wr_data_rom[  277]='h00000111;
    rd_cycle[  278] = 1'b1;  wr_cycle[  278] = 1'b0;  addr_rom[  278]='h00000060;  wr_data_rom[  278]='h00000000;
    rd_cycle[  279] = 1'b0;  wr_cycle[  279] = 1'b1;  addr_rom[  279]='h0000013c;  wr_data_rom[  279]='h000000f4;
    rd_cycle[  280] = 1'b1;  wr_cycle[  280] = 1'b0;  addr_rom[  280]='h0000005c;  wr_data_rom[  280]='h00000000;
    rd_cycle[  281] = 1'b0;  wr_cycle[  281] = 1'b1;  addr_rom[  281]='h0000003c;  wr_data_rom[  281]='h00000171;
    rd_cycle[  282] = 1'b0;  wr_cycle[  282] = 1'b1;  addr_rom[  282]='h00000018;  wr_data_rom[  282]='h00000135;
    rd_cycle[  283] = 1'b1;  wr_cycle[  283] = 1'b0;  addr_rom[  283]='h0000001c;  wr_data_rom[  283]='h00000000;
    rd_cycle[  284] = 1'b1;  wr_cycle[  284] = 1'b0;  addr_rom[  284]='h00000130;  wr_data_rom[  284]='h00000000;
    rd_cycle[  285] = 1'b0;  wr_cycle[  285] = 1'b1;  addr_rom[  285]='h0000017c;  wr_data_rom[  285]='h000000ad;
    rd_cycle[  286] = 1'b1;  wr_cycle[  286] = 1'b0;  addr_rom[  286]='h000000e0;  wr_data_rom[  286]='h00000000;
    rd_cycle[  287] = 1'b1;  wr_cycle[  287] = 1'b0;  addr_rom[  287]='h000000b0;  wr_data_rom[  287]='h00000000;
    rd_cycle[  288] = 1'b0;  wr_cycle[  288] = 1'b1;  addr_rom[  288]='h000000f0;  wr_data_rom[  288]='h0000002f;
    rd_cycle[  289] = 1'b1;  wr_cycle[  289] = 1'b0;  addr_rom[  289]='h000000dc;  wr_data_rom[  289]='h00000000;
    rd_cycle[  290] = 1'b1;  wr_cycle[  290] = 1'b0;  addr_rom[  290]='h00000160;  wr_data_rom[  290]='h00000000;
    rd_cycle[  291] = 1'b1;  wr_cycle[  291] = 1'b0;  addr_rom[  291]='h00000110;  wr_data_rom[  291]='h00000000;
    rd_cycle[  292] = 1'b0;  wr_cycle[  292] = 1'b1;  addr_rom[  292]='h000000dc;  wr_data_rom[  292]='h00000027;
    rd_cycle[  293] = 1'b0;  wr_cycle[  293] = 1'b1;  addr_rom[  293]='h00000104;  wr_data_rom[  293]='h0000015d;
    rd_cycle[  294] = 1'b0;  wr_cycle[  294] = 1'b1;  addr_rom[  294]='h000000b8;  wr_data_rom[  294]='h0000007b;
    rd_cycle[  295] = 1'b1;  wr_cycle[  295] = 1'b0;  addr_rom[  295]='h0000011c;  wr_data_rom[  295]='h00000000;
    rd_cycle[  296] = 1'b0;  wr_cycle[  296] = 1'b1;  addr_rom[  296]='h00000120;  wr_data_rom[  296]='h00000189;
    rd_cycle[  297] = 1'b1;  wr_cycle[  297] = 1'b0;  addr_rom[  297]='h00000154;  wr_data_rom[  297]='h00000000;
    rd_cycle[  298] = 1'b0;  wr_cycle[  298] = 1'b1;  addr_rom[  298]='h0000006c;  wr_data_rom[  298]='h0000004c;
    rd_cycle[  299] = 1'b0;  wr_cycle[  299] = 1'b1;  addr_rom[  299]='h000000c8;  wr_data_rom[  299]='h000000b2;
    rd_cycle[  300] = 1'b0;  wr_cycle[  300] = 1'b1;  addr_rom[  300]='h00000144;  wr_data_rom[  300]='h000000d5;
    rd_cycle[  301] = 1'b1;  wr_cycle[  301] = 1'b0;  addr_rom[  301]='h000000bc;  wr_data_rom[  301]='h00000000;
    rd_cycle[  302] = 1'b0;  wr_cycle[  302] = 1'b1;  addr_rom[  302]='h000000e4;  wr_data_rom[  302]='h0000006a;
    rd_cycle[  303] = 1'b0;  wr_cycle[  303] = 1'b1;  addr_rom[  303]='h000000e4;  wr_data_rom[  303]='h00000123;
    rd_cycle[  304] = 1'b0;  wr_cycle[  304] = 1'b1;  addr_rom[  304]='h0000000c;  wr_data_rom[  304]='h00000129;
    rd_cycle[  305] = 1'b1;  wr_cycle[  305] = 1'b0;  addr_rom[  305]='h00000008;  wr_data_rom[  305]='h00000000;
    rd_cycle[  306] = 1'b1;  wr_cycle[  306] = 1'b0;  addr_rom[  306]='h000000b8;  wr_data_rom[  306]='h00000000;
    rd_cycle[  307] = 1'b0;  wr_cycle[  307] = 1'b1;  addr_rom[  307]='h00000078;  wr_data_rom[  307]='h0000006c;
    rd_cycle[  308] = 1'b0;  wr_cycle[  308] = 1'b1;  addr_rom[  308]='h0000018c;  wr_data_rom[  308]='h0000004e;
    rd_cycle[  309] = 1'b0;  wr_cycle[  309] = 1'b1;  addr_rom[  309]='h0000016c;  wr_data_rom[  309]='h0000014f;
    rd_cycle[  310] = 1'b0;  wr_cycle[  310] = 1'b1;  addr_rom[  310]='h0000018c;  wr_data_rom[  310]='h0000008a;
    rd_cycle[  311] = 1'b1;  wr_cycle[  311] = 1'b0;  addr_rom[  311]='h00000080;  wr_data_rom[  311]='h00000000;
    rd_cycle[  312] = 1'b1;  wr_cycle[  312] = 1'b0;  addr_rom[  312]='h000000b8;  wr_data_rom[  312]='h00000000;
    rd_cycle[  313] = 1'b1;  wr_cycle[  313] = 1'b0;  addr_rom[  313]='h00000164;  wr_data_rom[  313]='h00000000;
    rd_cycle[  314] = 1'b0;  wr_cycle[  314] = 1'b1;  addr_rom[  314]='h000000c0;  wr_data_rom[  314]='h0000007f;
    rd_cycle[  315] = 1'b0;  wr_cycle[  315] = 1'b1;  addr_rom[  315]='h00000138;  wr_data_rom[  315]='h00000000;
    rd_cycle[  316] = 1'b1;  wr_cycle[  316] = 1'b0;  addr_rom[  316]='h00000048;  wr_data_rom[  316]='h00000000;
    rd_cycle[  317] = 1'b0;  wr_cycle[  317] = 1'b1;  addr_rom[  317]='h00000040;  wr_data_rom[  317]='h000000e9;
    rd_cycle[  318] = 1'b1;  wr_cycle[  318] = 1'b0;  addr_rom[  318]='h00000074;  wr_data_rom[  318]='h00000000;
    rd_cycle[  319] = 1'b0;  wr_cycle[  319] = 1'b1;  addr_rom[  319]='h0000004c;  wr_data_rom[  319]='h00000087;
    rd_cycle[  320] = 1'b0;  wr_cycle[  320] = 1'b1;  addr_rom[  320]='h00000184;  wr_data_rom[  320]='h00000171;
    rd_cycle[  321] = 1'b1;  wr_cycle[  321] = 1'b0;  addr_rom[  321]='h00000158;  wr_data_rom[  321]='h00000000;
    rd_cycle[  322] = 1'b0;  wr_cycle[  322] = 1'b1;  addr_rom[  322]='h000000f8;  wr_data_rom[  322]='h0000008f;
    rd_cycle[  323] = 1'b0;  wr_cycle[  323] = 1'b1;  addr_rom[  323]='h00000078;  wr_data_rom[  323]='h00000115;
    rd_cycle[  324] = 1'b1;  wr_cycle[  324] = 1'b0;  addr_rom[  324]='h0000015c;  wr_data_rom[  324]='h00000000;
    rd_cycle[  325] = 1'b0;  wr_cycle[  325] = 1'b1;  addr_rom[  325]='h00000060;  wr_data_rom[  325]='h00000057;
    rd_cycle[  326] = 1'b0;  wr_cycle[  326] = 1'b1;  addr_rom[  326]='h00000154;  wr_data_rom[  326]='h000000ef;
    rd_cycle[  327] = 1'b0;  wr_cycle[  327] = 1'b1;  addr_rom[  327]='h0000002c;  wr_data_rom[  327]='h000000c3;
    rd_cycle[  328] = 1'b0;  wr_cycle[  328] = 1'b1;  addr_rom[  328]='h00000020;  wr_data_rom[  328]='h000000a4;
    rd_cycle[  329] = 1'b1;  wr_cycle[  329] = 1'b0;  addr_rom[  329]='h00000038;  wr_data_rom[  329]='h00000000;
    rd_cycle[  330] = 1'b1;  wr_cycle[  330] = 1'b0;  addr_rom[  330]='h00000104;  wr_data_rom[  330]='h00000000;
    rd_cycle[  331] = 1'b1;  wr_cycle[  331] = 1'b0;  addr_rom[  331]='h00000138;  wr_data_rom[  331]='h00000000;
    rd_cycle[  332] = 1'b1;  wr_cycle[  332] = 1'b0;  addr_rom[  332]='h00000120;  wr_data_rom[  332]='h00000000;
    rd_cycle[  333] = 1'b1;  wr_cycle[  333] = 1'b0;  addr_rom[  333]='h00000140;  wr_data_rom[  333]='h00000000;
    rd_cycle[  334] = 1'b1;  wr_cycle[  334] = 1'b0;  addr_rom[  334]='h0000001c;  wr_data_rom[  334]='h00000000;
    rd_cycle[  335] = 1'b0;  wr_cycle[  335] = 1'b1;  addr_rom[  335]='h00000124;  wr_data_rom[  335]='h00000117;
    rd_cycle[  336] = 1'b0;  wr_cycle[  336] = 1'b1;  addr_rom[  336]='h000000cc;  wr_data_rom[  336]='h00000144;
    rd_cycle[  337] = 1'b0;  wr_cycle[  337] = 1'b1;  addr_rom[  337]='h0000015c;  wr_data_rom[  337]='h00000021;
    rd_cycle[  338] = 1'b0;  wr_cycle[  338] = 1'b1;  addr_rom[  338]='h00000134;  wr_data_rom[  338]='h00000138;
    rd_cycle[  339] = 1'b1;  wr_cycle[  339] = 1'b0;  addr_rom[  339]='h0000013c;  wr_data_rom[  339]='h00000000;
    rd_cycle[  340] = 1'b0;  wr_cycle[  340] = 1'b1;  addr_rom[  340]='h0000018c;  wr_data_rom[  340]='h00000122;
    rd_cycle[  341] = 1'b0;  wr_cycle[  341] = 1'b1;  addr_rom[  341]='h00000120;  wr_data_rom[  341]='h0000005d;
    rd_cycle[  342] = 1'b1;  wr_cycle[  342] = 1'b0;  addr_rom[  342]='h000000fc;  wr_data_rom[  342]='h00000000;
    rd_cycle[  343] = 1'b1;  wr_cycle[  343] = 1'b0;  addr_rom[  343]='h000000a4;  wr_data_rom[  343]='h00000000;
    rd_cycle[  344] = 1'b0;  wr_cycle[  344] = 1'b1;  addr_rom[  344]='h00000084;  wr_data_rom[  344]='h000000f9;
    rd_cycle[  345] = 1'b0;  wr_cycle[  345] = 1'b1;  addr_rom[  345]='h0000018c;  wr_data_rom[  345]='h00000009;
    rd_cycle[  346] = 1'b0;  wr_cycle[  346] = 1'b1;  addr_rom[  346]='h0000003c;  wr_data_rom[  346]='h0000011e;
    rd_cycle[  347] = 1'b1;  wr_cycle[  347] = 1'b0;  addr_rom[  347]='h00000118;  wr_data_rom[  347]='h00000000;
    rd_cycle[  348] = 1'b1;  wr_cycle[  348] = 1'b0;  addr_rom[  348]='h000000d0;  wr_data_rom[  348]='h00000000;
    rd_cycle[  349] = 1'b1;  wr_cycle[  349] = 1'b0;  addr_rom[  349]='h000000d8;  wr_data_rom[  349]='h00000000;
    rd_cycle[  350] = 1'b0;  wr_cycle[  350] = 1'b1;  addr_rom[  350]='h0000008c;  wr_data_rom[  350]='h00000059;
    rd_cycle[  351] = 1'b0;  wr_cycle[  351] = 1'b1;  addr_rom[  351]='h0000016c;  wr_data_rom[  351]='h000000e1;
    rd_cycle[  352] = 1'b0;  wr_cycle[  352] = 1'b1;  addr_rom[  352]='h00000188;  wr_data_rom[  352]='h0000005d;
    rd_cycle[  353] = 1'b1;  wr_cycle[  353] = 1'b0;  addr_rom[  353]='h00000048;  wr_data_rom[  353]='h00000000;
    rd_cycle[  354] = 1'b1;  wr_cycle[  354] = 1'b0;  addr_rom[  354]='h0000001c;  wr_data_rom[  354]='h00000000;
    rd_cycle[  355] = 1'b0;  wr_cycle[  355] = 1'b1;  addr_rom[  355]='h00000074;  wr_data_rom[  355]='h000000a3;
    rd_cycle[  356] = 1'b0;  wr_cycle[  356] = 1'b1;  addr_rom[  356]='h00000148;  wr_data_rom[  356]='h000000ba;
    rd_cycle[  357] = 1'b1;  wr_cycle[  357] = 1'b0;  addr_rom[  357]='h000000c4;  wr_data_rom[  357]='h00000000;
    rd_cycle[  358] = 1'b0;  wr_cycle[  358] = 1'b1;  addr_rom[  358]='h00000050;  wr_data_rom[  358]='h00000119;
    rd_cycle[  359] = 1'b1;  wr_cycle[  359] = 1'b0;  addr_rom[  359]='h000000f8;  wr_data_rom[  359]='h00000000;
    rd_cycle[  360] = 1'b1;  wr_cycle[  360] = 1'b0;  addr_rom[  360]='h00000004;  wr_data_rom[  360]='h00000000;
    rd_cycle[  361] = 1'b1;  wr_cycle[  361] = 1'b0;  addr_rom[  361]='h00000050;  wr_data_rom[  361]='h00000000;
    rd_cycle[  362] = 1'b0;  wr_cycle[  362] = 1'b1;  addr_rom[  362]='h00000160;  wr_data_rom[  362]='h00000013;
    rd_cycle[  363] = 1'b0;  wr_cycle[  363] = 1'b1;  addr_rom[  363]='h00000038;  wr_data_rom[  363]='h00000188;
    rd_cycle[  364] = 1'b0;  wr_cycle[  364] = 1'b1;  addr_rom[  364]='h000000e8;  wr_data_rom[  364]='h00000163;
    rd_cycle[  365] = 1'b0;  wr_cycle[  365] = 1'b1;  addr_rom[  365]='h00000090;  wr_data_rom[  365]='h00000067;
    rd_cycle[  366] = 1'b0;  wr_cycle[  366] = 1'b1;  addr_rom[  366]='h000000c8;  wr_data_rom[  366]='h0000001e;
    rd_cycle[  367] = 1'b0;  wr_cycle[  367] = 1'b1;  addr_rom[  367]='h0000001c;  wr_data_rom[  367]='h00000008;
    rd_cycle[  368] = 1'b1;  wr_cycle[  368] = 1'b0;  addr_rom[  368]='h00000094;  wr_data_rom[  368]='h00000000;
    rd_cycle[  369] = 1'b0;  wr_cycle[  369] = 1'b1;  addr_rom[  369]='h00000128;  wr_data_rom[  369]='h0000015f;
    rd_cycle[  370] = 1'b1;  wr_cycle[  370] = 1'b0;  addr_rom[  370]='h0000003c;  wr_data_rom[  370]='h00000000;
    rd_cycle[  371] = 1'b0;  wr_cycle[  371] = 1'b1;  addr_rom[  371]='h0000006c;  wr_data_rom[  371]='h000000ba;
    rd_cycle[  372] = 1'b0;  wr_cycle[  372] = 1'b1;  addr_rom[  372]='h00000068;  wr_data_rom[  372]='h0000008a;
    rd_cycle[  373] = 1'b0;  wr_cycle[  373] = 1'b1;  addr_rom[  373]='h000000a8;  wr_data_rom[  373]='h000000c1;
    rd_cycle[  374] = 1'b0;  wr_cycle[  374] = 1'b1;  addr_rom[  374]='h0000002c;  wr_data_rom[  374]='h00000075;
    rd_cycle[  375] = 1'b1;  wr_cycle[  375] = 1'b0;  addr_rom[  375]='h00000060;  wr_data_rom[  375]='h00000000;
    rd_cycle[  376] = 1'b0;  wr_cycle[  376] = 1'b1;  addr_rom[  376]='h00000004;  wr_data_rom[  376]='h000000ef;
    rd_cycle[  377] = 1'b1;  wr_cycle[  377] = 1'b0;  addr_rom[  377]='h00000080;  wr_data_rom[  377]='h00000000;
    rd_cycle[  378] = 1'b0;  wr_cycle[  378] = 1'b1;  addr_rom[  378]='h00000028;  wr_data_rom[  378]='h00000070;
    rd_cycle[  379] = 1'b0;  wr_cycle[  379] = 1'b1;  addr_rom[  379]='h000000b0;  wr_data_rom[  379]='h00000134;
    rd_cycle[  380] = 1'b1;  wr_cycle[  380] = 1'b0;  addr_rom[  380]='h00000070;  wr_data_rom[  380]='h00000000;
    rd_cycle[  381] = 1'b0;  wr_cycle[  381] = 1'b1;  addr_rom[  381]='h000000b8;  wr_data_rom[  381]='h00000136;
    rd_cycle[  382] = 1'b1;  wr_cycle[  382] = 1'b0;  addr_rom[  382]='h000000ac;  wr_data_rom[  382]='h00000000;
    rd_cycle[  383] = 1'b1;  wr_cycle[  383] = 1'b0;  addr_rom[  383]='h00000180;  wr_data_rom[  383]='h00000000;
    rd_cycle[  384] = 1'b0;  wr_cycle[  384] = 1'b1;  addr_rom[  384]='h00000104;  wr_data_rom[  384]='h00000146;
    rd_cycle[  385] = 1'b1;  wr_cycle[  385] = 1'b0;  addr_rom[  385]='h00000070;  wr_data_rom[  385]='h00000000;
    rd_cycle[  386] = 1'b0;  wr_cycle[  386] = 1'b1;  addr_rom[  386]='h000000f8;  wr_data_rom[  386]='h000000ad;
    rd_cycle[  387] = 1'b0;  wr_cycle[  387] = 1'b1;  addr_rom[  387]='h00000028;  wr_data_rom[  387]='h00000006;
    rd_cycle[  388] = 1'b1;  wr_cycle[  388] = 1'b0;  addr_rom[  388]='h00000134;  wr_data_rom[  388]='h00000000;
    rd_cycle[  389] = 1'b0;  wr_cycle[  389] = 1'b1;  addr_rom[  389]='h000000d4;  wr_data_rom[  389]='h0000014d;
    rd_cycle[  390] = 1'b0;  wr_cycle[  390] = 1'b1;  addr_rom[  390]='h00000054;  wr_data_rom[  390]='h0000002e;
    rd_cycle[  391] = 1'b1;  wr_cycle[  391] = 1'b0;  addr_rom[  391]='h00000078;  wr_data_rom[  391]='h00000000;
    rd_cycle[  392] = 1'b1;  wr_cycle[  392] = 1'b0;  addr_rom[  392]='h000000ac;  wr_data_rom[  392]='h00000000;
    rd_cycle[  393] = 1'b1;  wr_cycle[  393] = 1'b0;  addr_rom[  393]='h00000130;  wr_data_rom[  393]='h00000000;
    rd_cycle[  394] = 1'b1;  wr_cycle[  394] = 1'b0;  addr_rom[  394]='h00000028;  wr_data_rom[  394]='h00000000;
    rd_cycle[  395] = 1'b1;  wr_cycle[  395] = 1'b0;  addr_rom[  395]='h000000d8;  wr_data_rom[  395]='h00000000;
    rd_cycle[  396] = 1'b1;  wr_cycle[  396] = 1'b0;  addr_rom[  396]='h00000150;  wr_data_rom[  396]='h00000000;
    rd_cycle[  397] = 1'b1;  wr_cycle[  397] = 1'b0;  addr_rom[  397]='h00000118;  wr_data_rom[  397]='h00000000;
    rd_cycle[  398] = 1'b0;  wr_cycle[  398] = 1'b1;  addr_rom[  398]='h0000010c;  wr_data_rom[  398]='h000000b0;
    rd_cycle[  399] = 1'b1;  wr_cycle[  399] = 1'b0;  addr_rom[  399]='h00000048;  wr_data_rom[  399]='h00000000;
    // 100 silence cycles
    rd_cycle[  400] = 1'b0;  wr_cycle[  400] = 1'b0;  addr_rom[  400]='h00000000;  wr_data_rom[  400]='h00000000;
    rd_cycle[  401] = 1'b0;  wr_cycle[  401] = 1'b0;  addr_rom[  401]='h00000000;  wr_data_rom[  401]='h00000000;
    rd_cycle[  402] = 1'b0;  wr_cycle[  402] = 1'b0;  addr_rom[  402]='h00000000;  wr_data_rom[  402]='h00000000;
    rd_cycle[  403] = 1'b0;  wr_cycle[  403] = 1'b0;  addr_rom[  403]='h00000000;  wr_data_rom[  403]='h00000000;
    rd_cycle[  404] = 1'b0;  wr_cycle[  404] = 1'b0;  addr_rom[  404]='h00000000;  wr_data_rom[  404]='h00000000;
    rd_cycle[  405] = 1'b0;  wr_cycle[  405] = 1'b0;  addr_rom[  405]='h00000000;  wr_data_rom[  405]='h00000000;
    rd_cycle[  406] = 1'b0;  wr_cycle[  406] = 1'b0;  addr_rom[  406]='h00000000;  wr_data_rom[  406]='h00000000;
    rd_cycle[  407] = 1'b0;  wr_cycle[  407] = 1'b0;  addr_rom[  407]='h00000000;  wr_data_rom[  407]='h00000000;
    rd_cycle[  408] = 1'b0;  wr_cycle[  408] = 1'b0;  addr_rom[  408]='h00000000;  wr_data_rom[  408]='h00000000;
    rd_cycle[  409] = 1'b0;  wr_cycle[  409] = 1'b0;  addr_rom[  409]='h00000000;  wr_data_rom[  409]='h00000000;
    rd_cycle[  410] = 1'b0;  wr_cycle[  410] = 1'b0;  addr_rom[  410]='h00000000;  wr_data_rom[  410]='h00000000;
    rd_cycle[  411] = 1'b0;  wr_cycle[  411] = 1'b0;  addr_rom[  411]='h00000000;  wr_data_rom[  411]='h00000000;
    rd_cycle[  412] = 1'b0;  wr_cycle[  412] = 1'b0;  addr_rom[  412]='h00000000;  wr_data_rom[  412]='h00000000;
    rd_cycle[  413] = 1'b0;  wr_cycle[  413] = 1'b0;  addr_rom[  413]='h00000000;  wr_data_rom[  413]='h00000000;
    rd_cycle[  414] = 1'b0;  wr_cycle[  414] = 1'b0;  addr_rom[  414]='h00000000;  wr_data_rom[  414]='h00000000;
    rd_cycle[  415] = 1'b0;  wr_cycle[  415] = 1'b0;  addr_rom[  415]='h00000000;  wr_data_rom[  415]='h00000000;
    rd_cycle[  416] = 1'b0;  wr_cycle[  416] = 1'b0;  addr_rom[  416]='h00000000;  wr_data_rom[  416]='h00000000;
    rd_cycle[  417] = 1'b0;  wr_cycle[  417] = 1'b0;  addr_rom[  417]='h00000000;  wr_data_rom[  417]='h00000000;
    rd_cycle[  418] = 1'b0;  wr_cycle[  418] = 1'b0;  addr_rom[  418]='h00000000;  wr_data_rom[  418]='h00000000;
    rd_cycle[  419] = 1'b0;  wr_cycle[  419] = 1'b0;  addr_rom[  419]='h00000000;  wr_data_rom[  419]='h00000000;
    rd_cycle[  420] = 1'b0;  wr_cycle[  420] = 1'b0;  addr_rom[  420]='h00000000;  wr_data_rom[  420]='h00000000;
    rd_cycle[  421] = 1'b0;  wr_cycle[  421] = 1'b0;  addr_rom[  421]='h00000000;  wr_data_rom[  421]='h00000000;
    rd_cycle[  422] = 1'b0;  wr_cycle[  422] = 1'b0;  addr_rom[  422]='h00000000;  wr_data_rom[  422]='h00000000;
    rd_cycle[  423] = 1'b0;  wr_cycle[  423] = 1'b0;  addr_rom[  423]='h00000000;  wr_data_rom[  423]='h00000000;
    rd_cycle[  424] = 1'b0;  wr_cycle[  424] = 1'b0;  addr_rom[  424]='h00000000;  wr_data_rom[  424]='h00000000;
    rd_cycle[  425] = 1'b0;  wr_cycle[  425] = 1'b0;  addr_rom[  425]='h00000000;  wr_data_rom[  425]='h00000000;
    rd_cycle[  426] = 1'b0;  wr_cycle[  426] = 1'b0;  addr_rom[  426]='h00000000;  wr_data_rom[  426]='h00000000;
    rd_cycle[  427] = 1'b0;  wr_cycle[  427] = 1'b0;  addr_rom[  427]='h00000000;  wr_data_rom[  427]='h00000000;
    rd_cycle[  428] = 1'b0;  wr_cycle[  428] = 1'b0;  addr_rom[  428]='h00000000;  wr_data_rom[  428]='h00000000;
    rd_cycle[  429] = 1'b0;  wr_cycle[  429] = 1'b0;  addr_rom[  429]='h00000000;  wr_data_rom[  429]='h00000000;
    rd_cycle[  430] = 1'b0;  wr_cycle[  430] = 1'b0;  addr_rom[  430]='h00000000;  wr_data_rom[  430]='h00000000;
    rd_cycle[  431] = 1'b0;  wr_cycle[  431] = 1'b0;  addr_rom[  431]='h00000000;  wr_data_rom[  431]='h00000000;
    rd_cycle[  432] = 1'b0;  wr_cycle[  432] = 1'b0;  addr_rom[  432]='h00000000;  wr_data_rom[  432]='h00000000;
    rd_cycle[  433] = 1'b0;  wr_cycle[  433] = 1'b0;  addr_rom[  433]='h00000000;  wr_data_rom[  433]='h00000000;
    rd_cycle[  434] = 1'b0;  wr_cycle[  434] = 1'b0;  addr_rom[  434]='h00000000;  wr_data_rom[  434]='h00000000;
    rd_cycle[  435] = 1'b0;  wr_cycle[  435] = 1'b0;  addr_rom[  435]='h00000000;  wr_data_rom[  435]='h00000000;
    rd_cycle[  436] = 1'b0;  wr_cycle[  436] = 1'b0;  addr_rom[  436]='h00000000;  wr_data_rom[  436]='h00000000;
    rd_cycle[  437] = 1'b0;  wr_cycle[  437] = 1'b0;  addr_rom[  437]='h00000000;  wr_data_rom[  437]='h00000000;
    rd_cycle[  438] = 1'b0;  wr_cycle[  438] = 1'b0;  addr_rom[  438]='h00000000;  wr_data_rom[  438]='h00000000;
    rd_cycle[  439] = 1'b0;  wr_cycle[  439] = 1'b0;  addr_rom[  439]='h00000000;  wr_data_rom[  439]='h00000000;
    rd_cycle[  440] = 1'b0;  wr_cycle[  440] = 1'b0;  addr_rom[  440]='h00000000;  wr_data_rom[  440]='h00000000;
    rd_cycle[  441] = 1'b0;  wr_cycle[  441] = 1'b0;  addr_rom[  441]='h00000000;  wr_data_rom[  441]='h00000000;
    rd_cycle[  442] = 1'b0;  wr_cycle[  442] = 1'b0;  addr_rom[  442]='h00000000;  wr_data_rom[  442]='h00000000;
    rd_cycle[  443] = 1'b0;  wr_cycle[  443] = 1'b0;  addr_rom[  443]='h00000000;  wr_data_rom[  443]='h00000000;
    rd_cycle[  444] = 1'b0;  wr_cycle[  444] = 1'b0;  addr_rom[  444]='h00000000;  wr_data_rom[  444]='h00000000;
    rd_cycle[  445] = 1'b0;  wr_cycle[  445] = 1'b0;  addr_rom[  445]='h00000000;  wr_data_rom[  445]='h00000000;
    rd_cycle[  446] = 1'b0;  wr_cycle[  446] = 1'b0;  addr_rom[  446]='h00000000;  wr_data_rom[  446]='h00000000;
    rd_cycle[  447] = 1'b0;  wr_cycle[  447] = 1'b0;  addr_rom[  447]='h00000000;  wr_data_rom[  447]='h00000000;
    rd_cycle[  448] = 1'b0;  wr_cycle[  448] = 1'b0;  addr_rom[  448]='h00000000;  wr_data_rom[  448]='h00000000;
    rd_cycle[  449] = 1'b0;  wr_cycle[  449] = 1'b0;  addr_rom[  449]='h00000000;  wr_data_rom[  449]='h00000000;
    rd_cycle[  450] = 1'b0;  wr_cycle[  450] = 1'b0;  addr_rom[  450]='h00000000;  wr_data_rom[  450]='h00000000;
    rd_cycle[  451] = 1'b0;  wr_cycle[  451] = 1'b0;  addr_rom[  451]='h00000000;  wr_data_rom[  451]='h00000000;
    rd_cycle[  452] = 1'b0;  wr_cycle[  452] = 1'b0;  addr_rom[  452]='h00000000;  wr_data_rom[  452]='h00000000;
    rd_cycle[  453] = 1'b0;  wr_cycle[  453] = 1'b0;  addr_rom[  453]='h00000000;  wr_data_rom[  453]='h00000000;
    rd_cycle[  454] = 1'b0;  wr_cycle[  454] = 1'b0;  addr_rom[  454]='h00000000;  wr_data_rom[  454]='h00000000;
    rd_cycle[  455] = 1'b0;  wr_cycle[  455] = 1'b0;  addr_rom[  455]='h00000000;  wr_data_rom[  455]='h00000000;
    rd_cycle[  456] = 1'b0;  wr_cycle[  456] = 1'b0;  addr_rom[  456]='h00000000;  wr_data_rom[  456]='h00000000;
    rd_cycle[  457] = 1'b0;  wr_cycle[  457] = 1'b0;  addr_rom[  457]='h00000000;  wr_data_rom[  457]='h00000000;
    rd_cycle[  458] = 1'b0;  wr_cycle[  458] = 1'b0;  addr_rom[  458]='h00000000;  wr_data_rom[  458]='h00000000;
    rd_cycle[  459] = 1'b0;  wr_cycle[  459] = 1'b0;  addr_rom[  459]='h00000000;  wr_data_rom[  459]='h00000000;
    rd_cycle[  460] = 1'b0;  wr_cycle[  460] = 1'b0;  addr_rom[  460]='h00000000;  wr_data_rom[  460]='h00000000;
    rd_cycle[  461] = 1'b0;  wr_cycle[  461] = 1'b0;  addr_rom[  461]='h00000000;  wr_data_rom[  461]='h00000000;
    rd_cycle[  462] = 1'b0;  wr_cycle[  462] = 1'b0;  addr_rom[  462]='h00000000;  wr_data_rom[  462]='h00000000;
    rd_cycle[  463] = 1'b0;  wr_cycle[  463] = 1'b0;  addr_rom[  463]='h00000000;  wr_data_rom[  463]='h00000000;
    rd_cycle[  464] = 1'b0;  wr_cycle[  464] = 1'b0;  addr_rom[  464]='h00000000;  wr_data_rom[  464]='h00000000;
    rd_cycle[  465] = 1'b0;  wr_cycle[  465] = 1'b0;  addr_rom[  465]='h00000000;  wr_data_rom[  465]='h00000000;
    rd_cycle[  466] = 1'b0;  wr_cycle[  466] = 1'b0;  addr_rom[  466]='h00000000;  wr_data_rom[  466]='h00000000;
    rd_cycle[  467] = 1'b0;  wr_cycle[  467] = 1'b0;  addr_rom[  467]='h00000000;  wr_data_rom[  467]='h00000000;
    rd_cycle[  468] = 1'b0;  wr_cycle[  468] = 1'b0;  addr_rom[  468]='h00000000;  wr_data_rom[  468]='h00000000;
    rd_cycle[  469] = 1'b0;  wr_cycle[  469] = 1'b0;  addr_rom[  469]='h00000000;  wr_data_rom[  469]='h00000000;
    rd_cycle[  470] = 1'b0;  wr_cycle[  470] = 1'b0;  addr_rom[  470]='h00000000;  wr_data_rom[  470]='h00000000;
    rd_cycle[  471] = 1'b0;  wr_cycle[  471] = 1'b0;  addr_rom[  471]='h00000000;  wr_data_rom[  471]='h00000000;
    rd_cycle[  472] = 1'b0;  wr_cycle[  472] = 1'b0;  addr_rom[  472]='h00000000;  wr_data_rom[  472]='h00000000;
    rd_cycle[  473] = 1'b0;  wr_cycle[  473] = 1'b0;  addr_rom[  473]='h00000000;  wr_data_rom[  473]='h00000000;
    rd_cycle[  474] = 1'b0;  wr_cycle[  474] = 1'b0;  addr_rom[  474]='h00000000;  wr_data_rom[  474]='h00000000;
    rd_cycle[  475] = 1'b0;  wr_cycle[  475] = 1'b0;  addr_rom[  475]='h00000000;  wr_data_rom[  475]='h00000000;
    rd_cycle[  476] = 1'b0;  wr_cycle[  476] = 1'b0;  addr_rom[  476]='h00000000;  wr_data_rom[  476]='h00000000;
    rd_cycle[  477] = 1'b0;  wr_cycle[  477] = 1'b0;  addr_rom[  477]='h00000000;  wr_data_rom[  477]='h00000000;
    rd_cycle[  478] = 1'b0;  wr_cycle[  478] = 1'b0;  addr_rom[  478]='h00000000;  wr_data_rom[  478]='h00000000;
    rd_cycle[  479] = 1'b0;  wr_cycle[  479] = 1'b0;  addr_rom[  479]='h00000000;  wr_data_rom[  479]='h00000000;
    rd_cycle[  480] = 1'b0;  wr_cycle[  480] = 1'b0;  addr_rom[  480]='h00000000;  wr_data_rom[  480]='h00000000;
    rd_cycle[  481] = 1'b0;  wr_cycle[  481] = 1'b0;  addr_rom[  481]='h00000000;  wr_data_rom[  481]='h00000000;
    rd_cycle[  482] = 1'b0;  wr_cycle[  482] = 1'b0;  addr_rom[  482]='h00000000;  wr_data_rom[  482]='h00000000;
    rd_cycle[  483] = 1'b0;  wr_cycle[  483] = 1'b0;  addr_rom[  483]='h00000000;  wr_data_rom[  483]='h00000000;
    rd_cycle[  484] = 1'b0;  wr_cycle[  484] = 1'b0;  addr_rom[  484]='h00000000;  wr_data_rom[  484]='h00000000;
    rd_cycle[  485] = 1'b0;  wr_cycle[  485] = 1'b0;  addr_rom[  485]='h00000000;  wr_data_rom[  485]='h00000000;
    rd_cycle[  486] = 1'b0;  wr_cycle[  486] = 1'b0;  addr_rom[  486]='h00000000;  wr_data_rom[  486]='h00000000;
    rd_cycle[  487] = 1'b0;  wr_cycle[  487] = 1'b0;  addr_rom[  487]='h00000000;  wr_data_rom[  487]='h00000000;
    rd_cycle[  488] = 1'b0;  wr_cycle[  488] = 1'b0;  addr_rom[  488]='h00000000;  wr_data_rom[  488]='h00000000;
    rd_cycle[  489] = 1'b0;  wr_cycle[  489] = 1'b0;  addr_rom[  489]='h00000000;  wr_data_rom[  489]='h00000000;
    rd_cycle[  490] = 1'b0;  wr_cycle[  490] = 1'b0;  addr_rom[  490]='h00000000;  wr_data_rom[  490]='h00000000;
    rd_cycle[  491] = 1'b0;  wr_cycle[  491] = 1'b0;  addr_rom[  491]='h00000000;  wr_data_rom[  491]='h00000000;
    rd_cycle[  492] = 1'b0;  wr_cycle[  492] = 1'b0;  addr_rom[  492]='h00000000;  wr_data_rom[  492]='h00000000;
    rd_cycle[  493] = 1'b0;  wr_cycle[  493] = 1'b0;  addr_rom[  493]='h00000000;  wr_data_rom[  493]='h00000000;
    rd_cycle[  494] = 1'b0;  wr_cycle[  494] = 1'b0;  addr_rom[  494]='h00000000;  wr_data_rom[  494]='h00000000;
    rd_cycle[  495] = 1'b0;  wr_cycle[  495] = 1'b0;  addr_rom[  495]='h00000000;  wr_data_rom[  495]='h00000000;
    rd_cycle[  496] = 1'b0;  wr_cycle[  496] = 1'b0;  addr_rom[  496]='h00000000;  wr_data_rom[  496]='h00000000;
    rd_cycle[  497] = 1'b0;  wr_cycle[  497] = 1'b0;  addr_rom[  497]='h00000000;  wr_data_rom[  497]='h00000000;
    rd_cycle[  498] = 1'b0;  wr_cycle[  498] = 1'b0;  addr_rom[  498]='h00000000;  wr_data_rom[  498]='h00000000;
    rd_cycle[  499] = 1'b0;  wr_cycle[  499] = 1'b0;  addr_rom[  499]='h00000000;  wr_data_rom[  499]='h00000000;
    // 100 sequence read cycles
    rd_cycle[  500] = 1'b1;  wr_cycle[  500] = 1'b0;  addr_rom[  500]='h00000000;  wr_data_rom[  500]='h00000000;
    rd_cycle[  501] = 1'b1;  wr_cycle[  501] = 1'b0;  addr_rom[  501]='h00000004;  wr_data_rom[  501]='h00000000;
    rd_cycle[  502] = 1'b1;  wr_cycle[  502] = 1'b0;  addr_rom[  502]='h00000008;  wr_data_rom[  502]='h00000000;
    rd_cycle[  503] = 1'b1;  wr_cycle[  503] = 1'b0;  addr_rom[  503]='h0000000c;  wr_data_rom[  503]='h00000000;
    rd_cycle[  504] = 1'b1;  wr_cycle[  504] = 1'b0;  addr_rom[  504]='h00000010;  wr_data_rom[  504]='h00000000;
    rd_cycle[  505] = 1'b1;  wr_cycle[  505] = 1'b0;  addr_rom[  505]='h00000014;  wr_data_rom[  505]='h00000000;
    rd_cycle[  506] = 1'b1;  wr_cycle[  506] = 1'b0;  addr_rom[  506]='h00000018;  wr_data_rom[  506]='h00000000;
    rd_cycle[  507] = 1'b1;  wr_cycle[  507] = 1'b0;  addr_rom[  507]='h0000001c;  wr_data_rom[  507]='h00000000;
    rd_cycle[  508] = 1'b1;  wr_cycle[  508] = 1'b0;  addr_rom[  508]='h00000020;  wr_data_rom[  508]='h00000000;
    rd_cycle[  509] = 1'b1;  wr_cycle[  509] = 1'b0;  addr_rom[  509]='h00000024;  wr_data_rom[  509]='h00000000;
    rd_cycle[  510] = 1'b1;  wr_cycle[  510] = 1'b0;  addr_rom[  510]='h00000028;  wr_data_rom[  510]='h00000000;
    rd_cycle[  511] = 1'b1;  wr_cycle[  511] = 1'b0;  addr_rom[  511]='h0000002c;  wr_data_rom[  511]='h00000000;
    rd_cycle[  512] = 1'b1;  wr_cycle[  512] = 1'b0;  addr_rom[  512]='h00000030;  wr_data_rom[  512]='h00000000;
    rd_cycle[  513] = 1'b1;  wr_cycle[  513] = 1'b0;  addr_rom[  513]='h00000034;  wr_data_rom[  513]='h00000000;
    rd_cycle[  514] = 1'b1;  wr_cycle[  514] = 1'b0;  addr_rom[  514]='h00000038;  wr_data_rom[  514]='h00000000;
    rd_cycle[  515] = 1'b1;  wr_cycle[  515] = 1'b0;  addr_rom[  515]='h0000003c;  wr_data_rom[  515]='h00000000;
    rd_cycle[  516] = 1'b1;  wr_cycle[  516] = 1'b0;  addr_rom[  516]='h00000040;  wr_data_rom[  516]='h00000000;
    rd_cycle[  517] = 1'b1;  wr_cycle[  517] = 1'b0;  addr_rom[  517]='h00000044;  wr_data_rom[  517]='h00000000;
    rd_cycle[  518] = 1'b1;  wr_cycle[  518] = 1'b0;  addr_rom[  518]='h00000048;  wr_data_rom[  518]='h00000000;
    rd_cycle[  519] = 1'b1;  wr_cycle[  519] = 1'b0;  addr_rom[  519]='h0000004c;  wr_data_rom[  519]='h00000000;
    rd_cycle[  520] = 1'b1;  wr_cycle[  520] = 1'b0;  addr_rom[  520]='h00000050;  wr_data_rom[  520]='h00000000;
    rd_cycle[  521] = 1'b1;  wr_cycle[  521] = 1'b0;  addr_rom[  521]='h00000054;  wr_data_rom[  521]='h00000000;
    rd_cycle[  522] = 1'b1;  wr_cycle[  522] = 1'b0;  addr_rom[  522]='h00000058;  wr_data_rom[  522]='h00000000;
    rd_cycle[  523] = 1'b1;  wr_cycle[  523] = 1'b0;  addr_rom[  523]='h0000005c;  wr_data_rom[  523]='h00000000;
    rd_cycle[  524] = 1'b1;  wr_cycle[  524] = 1'b0;  addr_rom[  524]='h00000060;  wr_data_rom[  524]='h00000000;
    rd_cycle[  525] = 1'b1;  wr_cycle[  525] = 1'b0;  addr_rom[  525]='h00000064;  wr_data_rom[  525]='h00000000;
    rd_cycle[  526] = 1'b1;  wr_cycle[  526] = 1'b0;  addr_rom[  526]='h00000068;  wr_data_rom[  526]='h00000000;
    rd_cycle[  527] = 1'b1;  wr_cycle[  527] = 1'b0;  addr_rom[  527]='h0000006c;  wr_data_rom[  527]='h00000000;
    rd_cycle[  528] = 1'b1;  wr_cycle[  528] = 1'b0;  addr_rom[  528]='h00000070;  wr_data_rom[  528]='h00000000;
    rd_cycle[  529] = 1'b1;  wr_cycle[  529] = 1'b0;  addr_rom[  529]='h00000074;  wr_data_rom[  529]='h00000000;
    rd_cycle[  530] = 1'b1;  wr_cycle[  530] = 1'b0;  addr_rom[  530]='h00000078;  wr_data_rom[  530]='h00000000;
    rd_cycle[  531] = 1'b1;  wr_cycle[  531] = 1'b0;  addr_rom[  531]='h0000007c;  wr_data_rom[  531]='h00000000;
    rd_cycle[  532] = 1'b1;  wr_cycle[  532] = 1'b0;  addr_rom[  532]='h00000080;  wr_data_rom[  532]='h00000000;
    rd_cycle[  533] = 1'b1;  wr_cycle[  533] = 1'b0;  addr_rom[  533]='h00000084;  wr_data_rom[  533]='h00000000;
    rd_cycle[  534] = 1'b1;  wr_cycle[  534] = 1'b0;  addr_rom[  534]='h00000088;  wr_data_rom[  534]='h00000000;
    rd_cycle[  535] = 1'b1;  wr_cycle[  535] = 1'b0;  addr_rom[  535]='h0000008c;  wr_data_rom[  535]='h00000000;
    rd_cycle[  536] = 1'b1;  wr_cycle[  536] = 1'b0;  addr_rom[  536]='h00000090;  wr_data_rom[  536]='h00000000;
    rd_cycle[  537] = 1'b1;  wr_cycle[  537] = 1'b0;  addr_rom[  537]='h00000094;  wr_data_rom[  537]='h00000000;
    rd_cycle[  538] = 1'b1;  wr_cycle[  538] = 1'b0;  addr_rom[  538]='h00000098;  wr_data_rom[  538]='h00000000;
    rd_cycle[  539] = 1'b1;  wr_cycle[  539] = 1'b0;  addr_rom[  539]='h0000009c;  wr_data_rom[  539]='h00000000;
    rd_cycle[  540] = 1'b1;  wr_cycle[  540] = 1'b0;  addr_rom[  540]='h000000a0;  wr_data_rom[  540]='h00000000;
    rd_cycle[  541] = 1'b1;  wr_cycle[  541] = 1'b0;  addr_rom[  541]='h000000a4;  wr_data_rom[  541]='h00000000;
    rd_cycle[  542] = 1'b1;  wr_cycle[  542] = 1'b0;  addr_rom[  542]='h000000a8;  wr_data_rom[  542]='h00000000;
    rd_cycle[  543] = 1'b1;  wr_cycle[  543] = 1'b0;  addr_rom[  543]='h000000ac;  wr_data_rom[  543]='h00000000;
    rd_cycle[  544] = 1'b1;  wr_cycle[  544] = 1'b0;  addr_rom[  544]='h000000b0;  wr_data_rom[  544]='h00000000;
    rd_cycle[  545] = 1'b1;  wr_cycle[  545] = 1'b0;  addr_rom[  545]='h000000b4;  wr_data_rom[  545]='h00000000;
    rd_cycle[  546] = 1'b1;  wr_cycle[  546] = 1'b0;  addr_rom[  546]='h000000b8;  wr_data_rom[  546]='h00000000;
    rd_cycle[  547] = 1'b1;  wr_cycle[  547] = 1'b0;  addr_rom[  547]='h000000bc;  wr_data_rom[  547]='h00000000;
    rd_cycle[  548] = 1'b1;  wr_cycle[  548] = 1'b0;  addr_rom[  548]='h000000c0;  wr_data_rom[  548]='h00000000;
    rd_cycle[  549] = 1'b1;  wr_cycle[  549] = 1'b0;  addr_rom[  549]='h000000c4;  wr_data_rom[  549]='h00000000;
    rd_cycle[  550] = 1'b1;  wr_cycle[  550] = 1'b0;  addr_rom[  550]='h000000c8;  wr_data_rom[  550]='h00000000;
    rd_cycle[  551] = 1'b1;  wr_cycle[  551] = 1'b0;  addr_rom[  551]='h000000cc;  wr_data_rom[  551]='h00000000;
    rd_cycle[  552] = 1'b1;  wr_cycle[  552] = 1'b0;  addr_rom[  552]='h000000d0;  wr_data_rom[  552]='h00000000;
    rd_cycle[  553] = 1'b1;  wr_cycle[  553] = 1'b0;  addr_rom[  553]='h000000d4;  wr_data_rom[  553]='h00000000;
    rd_cycle[  554] = 1'b1;  wr_cycle[  554] = 1'b0;  addr_rom[  554]='h000000d8;  wr_data_rom[  554]='h00000000;
    rd_cycle[  555] = 1'b1;  wr_cycle[  555] = 1'b0;  addr_rom[  555]='h000000dc;  wr_data_rom[  555]='h00000000;
    rd_cycle[  556] = 1'b1;  wr_cycle[  556] = 1'b0;  addr_rom[  556]='h000000e0;  wr_data_rom[  556]='h00000000;
    rd_cycle[  557] = 1'b1;  wr_cycle[  557] = 1'b0;  addr_rom[  557]='h000000e4;  wr_data_rom[  557]='h00000000;
    rd_cycle[  558] = 1'b1;  wr_cycle[  558] = 1'b0;  addr_rom[  558]='h000000e8;  wr_data_rom[  558]='h00000000;
    rd_cycle[  559] = 1'b1;  wr_cycle[  559] = 1'b0;  addr_rom[  559]='h000000ec;  wr_data_rom[  559]='h00000000;
    rd_cycle[  560] = 1'b1;  wr_cycle[  560] = 1'b0;  addr_rom[  560]='h000000f0;  wr_data_rom[  560]='h00000000;
    rd_cycle[  561] = 1'b1;  wr_cycle[  561] = 1'b0;  addr_rom[  561]='h000000f4;  wr_data_rom[  561]='h00000000;
    rd_cycle[  562] = 1'b1;  wr_cycle[  562] = 1'b0;  addr_rom[  562]='h000000f8;  wr_data_rom[  562]='h00000000;
    rd_cycle[  563] = 1'b1;  wr_cycle[  563] = 1'b0;  addr_rom[  563]='h000000fc;  wr_data_rom[  563]='h00000000;
    rd_cycle[  564] = 1'b1;  wr_cycle[  564] = 1'b0;  addr_rom[  564]='h00000100;  wr_data_rom[  564]='h00000000;
    rd_cycle[  565] = 1'b1;  wr_cycle[  565] = 1'b0;  addr_rom[  565]='h00000104;  wr_data_rom[  565]='h00000000;
    rd_cycle[  566] = 1'b1;  wr_cycle[  566] = 1'b0;  addr_rom[  566]='h00000108;  wr_data_rom[  566]='h00000000;
    rd_cycle[  567] = 1'b1;  wr_cycle[  567] = 1'b0;  addr_rom[  567]='h0000010c;  wr_data_rom[  567]='h00000000;
    rd_cycle[  568] = 1'b1;  wr_cycle[  568] = 1'b0;  addr_rom[  568]='h00000110;  wr_data_rom[  568]='h00000000;
    rd_cycle[  569] = 1'b1;  wr_cycle[  569] = 1'b0;  addr_rom[  569]='h00000114;  wr_data_rom[  569]='h00000000;
    rd_cycle[  570] = 1'b1;  wr_cycle[  570] = 1'b0;  addr_rom[  570]='h00000118;  wr_data_rom[  570]='h00000000;
    rd_cycle[  571] = 1'b1;  wr_cycle[  571] = 1'b0;  addr_rom[  571]='h0000011c;  wr_data_rom[  571]='h00000000;
    rd_cycle[  572] = 1'b1;  wr_cycle[  572] = 1'b0;  addr_rom[  572]='h00000120;  wr_data_rom[  572]='h00000000;
    rd_cycle[  573] = 1'b1;  wr_cycle[  573] = 1'b0;  addr_rom[  573]='h00000124;  wr_data_rom[  573]='h00000000;
    rd_cycle[  574] = 1'b1;  wr_cycle[  574] = 1'b0;  addr_rom[  574]='h00000128;  wr_data_rom[  574]='h00000000;
    rd_cycle[  575] = 1'b1;  wr_cycle[  575] = 1'b0;  addr_rom[  575]='h0000012c;  wr_data_rom[  575]='h00000000;
    rd_cycle[  576] = 1'b1;  wr_cycle[  576] = 1'b0;  addr_rom[  576]='h00000130;  wr_data_rom[  576]='h00000000;
    rd_cycle[  577] = 1'b1;  wr_cycle[  577] = 1'b0;  addr_rom[  577]='h00000134;  wr_data_rom[  577]='h00000000;
    rd_cycle[  578] = 1'b1;  wr_cycle[  578] = 1'b0;  addr_rom[  578]='h00000138;  wr_data_rom[  578]='h00000000;
    rd_cycle[  579] = 1'b1;  wr_cycle[  579] = 1'b0;  addr_rom[  579]='h0000013c;  wr_data_rom[  579]='h00000000;
    rd_cycle[  580] = 1'b1;  wr_cycle[  580] = 1'b0;  addr_rom[  580]='h00000140;  wr_data_rom[  580]='h00000000;
    rd_cycle[  581] = 1'b1;  wr_cycle[  581] = 1'b0;  addr_rom[  581]='h00000144;  wr_data_rom[  581]='h00000000;
    rd_cycle[  582] = 1'b1;  wr_cycle[  582] = 1'b0;  addr_rom[  582]='h00000148;  wr_data_rom[  582]='h00000000;
    rd_cycle[  583] = 1'b1;  wr_cycle[  583] = 1'b0;  addr_rom[  583]='h0000014c;  wr_data_rom[  583]='h00000000;
    rd_cycle[  584] = 1'b1;  wr_cycle[  584] = 1'b0;  addr_rom[  584]='h00000150;  wr_data_rom[  584]='h00000000;
    rd_cycle[  585] = 1'b1;  wr_cycle[  585] = 1'b0;  addr_rom[  585]='h00000154;  wr_data_rom[  585]='h00000000;
    rd_cycle[  586] = 1'b1;  wr_cycle[  586] = 1'b0;  addr_rom[  586]='h00000158;  wr_data_rom[  586]='h00000000;
    rd_cycle[  587] = 1'b1;  wr_cycle[  587] = 1'b0;  addr_rom[  587]='h0000015c;  wr_data_rom[  587]='h00000000;
    rd_cycle[  588] = 1'b1;  wr_cycle[  588] = 1'b0;  addr_rom[  588]='h00000160;  wr_data_rom[  588]='h00000000;
    rd_cycle[  589] = 1'b1;  wr_cycle[  589] = 1'b0;  addr_rom[  589]='h00000164;  wr_data_rom[  589]='h00000000;
    rd_cycle[  590] = 1'b1;  wr_cycle[  590] = 1'b0;  addr_rom[  590]='h00000168;  wr_data_rom[  590]='h00000000;
    rd_cycle[  591] = 1'b1;  wr_cycle[  591] = 1'b0;  addr_rom[  591]='h0000016c;  wr_data_rom[  591]='h00000000;
    rd_cycle[  592] = 1'b1;  wr_cycle[  592] = 1'b0;  addr_rom[  592]='h00000170;  wr_data_rom[  592]='h00000000;
    rd_cycle[  593] = 1'b1;  wr_cycle[  593] = 1'b0;  addr_rom[  593]='h00000174;  wr_data_rom[  593]='h00000000;
    rd_cycle[  594] = 1'b1;  wr_cycle[  594] = 1'b0;  addr_rom[  594]='h00000178;  wr_data_rom[  594]='h00000000;
    rd_cycle[  595] = 1'b1;  wr_cycle[  595] = 1'b0;  addr_rom[  595]='h0000017c;  wr_data_rom[  595]='h00000000;
    rd_cycle[  596] = 1'b1;  wr_cycle[  596] = 1'b0;  addr_rom[  596]='h00000180;  wr_data_rom[  596]='h00000000;
    rd_cycle[  597] = 1'b1;  wr_cycle[  597] = 1'b0;  addr_rom[  597]='h00000184;  wr_data_rom[  597]='h00000000;
    rd_cycle[  598] = 1'b1;  wr_cycle[  598] = 1'b0;  addr_rom[  598]='h00000188;  wr_data_rom[  598]='h00000000;
    rd_cycle[  599] = 1'b1;  wr_cycle[  599] = 1'b0;  addr_rom[  599]='h0000018c;  wr_data_rom[  599]='h00000000;
end

initial begin
    validation_data[    0] = 'h00000000; 
    validation_data[    1] = 'h000000ef; 
    validation_data[    2] = 'h00000048; 
    validation_data[    3] = 'h00000129; 
    validation_data[    4] = 'h000000e3; 
    validation_data[    5] = 'h0000012e; 
    validation_data[    6] = 'h00000135; 
    validation_data[    7] = 'h00000008; 
    validation_data[    8] = 'h000000a4; 
    validation_data[    9] = 'h00000068; 
    validation_data[   10] = 'h00000006; 
    validation_data[   11] = 'h00000075; 
    validation_data[   12] = 'h00000147; 
    validation_data[   13] = 'h000000a7; 
    validation_data[   14] = 'h00000188; 
    validation_data[   15] = 'h0000011e; 
    validation_data[   16] = 'h000000e9; 
    validation_data[   17] = 'h0000009d; 
    validation_data[   18] = 'h00000065; 
    validation_data[   19] = 'h00000087; 
    validation_data[   20] = 'h00000119; 
    validation_data[   21] = 'h0000002e; 
    validation_data[   22] = 'h00000010; 
    validation_data[   23] = 'h000000fe; 
    validation_data[   24] = 'h00000057; 
    validation_data[   25] = 'h00000161; 
    validation_data[   26] = 'h0000008a; 
    validation_data[   27] = 'h000000ba; 
    validation_data[   28] = 'h0000002e; 
    validation_data[   29] = 'h000000a3; 
    validation_data[   30] = 'h00000115; 
    validation_data[   31] = 'h00000127; 
    validation_data[   32] = 'h0000016e; 
    validation_data[   33] = 'h000000f9; 
    validation_data[   34] = 'h0000001c; 
    validation_data[   35] = 'h00000059; 
    validation_data[   36] = 'h00000067; 
    validation_data[   37] = 'h0000011e; 
    validation_data[   38] = 'h00000036; 
    validation_data[   39] = 'h00000098; 
    validation_data[   40] = 'h0000005f; 
    validation_data[   41] = 'h0000015d; 
    validation_data[   42] = 'h000000c1; 
    validation_data[   43] = 'h0000014d; 
    validation_data[   44] = 'h00000134; 
    validation_data[   45] = 'h000000ff; 
    validation_data[   46] = 'h00000136; 
    validation_data[   47] = 'h00000173; 
    validation_data[   48] = 'h0000007f; 
    validation_data[   49] = 'h0000003e; 
    validation_data[   50] = 'h0000001e; 
    validation_data[   51] = 'h00000144; 
    validation_data[   52] = 'h000000b0; 
    validation_data[   53] = 'h0000014d; 
    validation_data[   54] = 'h00000111; 
    validation_data[   55] = 'h00000027; 
    validation_data[   56] = 'h000000f9; 
    validation_data[   57] = 'h00000123; 
    validation_data[   58] = 'h00000163; 
    validation_data[   59] = 'h00000046; 
    validation_data[   60] = 'h0000002f; 
    validation_data[   61] = 'h0000013f; 
    validation_data[   62] = 'h000000ad; 
    validation_data[   63] = 'h0000001d; 
    validation_data[   64] = 'h0000015e; 
    validation_data[   65] = 'h00000146; 
    validation_data[   66] = 'h00000054; 
    validation_data[   67] = 'h000000b0; 
    validation_data[   68] = 'h0000015e; 
    validation_data[   69] = 'h000000fa; 
    validation_data[   70] = 'h00000173; 
    validation_data[   71] = 'h0000008b; 
    validation_data[   72] = 'h0000005d; 
    validation_data[   73] = 'h00000117; 
    validation_data[   74] = 'h0000015f; 
    validation_data[   75] = 'h000000aa; 
    validation_data[   76] = 'h00000156; 
    validation_data[   77] = 'h00000138; 
    validation_data[   78] = 'h00000000; 
    validation_data[   79] = 'h000000f4; 
    validation_data[   80] = 'h00000142; 
    validation_data[   81] = 'h000000d5; 
    validation_data[   82] = 'h000000ba; 
    validation_data[   83] = 'h00000056; 
    validation_data[   84] = 'h000000f9; 
    validation_data[   85] = 'h000000ef; 
    validation_data[   86] = 'h00000022; 
    validation_data[   87] = 'h00000021; 
    validation_data[   88] = 'h00000013; 
    validation_data[   89] = 'h000000bf; 
    validation_data[   90] = 'h00000091; 
    validation_data[   91] = 'h000000e1; 
    validation_data[   92] = 'h0000014d; 
    validation_data[   93] = 'h0000001b; 
    validation_data[   94] = 'h00000085; 
    validation_data[   95] = 'h000000ad; 
    validation_data[   96] = 'h000000c1; 
    validation_data[   97] = 'h00000171; 
    validation_data[   98] = 'h0000005d; 
    validation_data[   99] = 'h00000009; 

end


reg clk = 1'b1, rst = 1'b1;
initial #4 rst = 1'b0;
always  #1 clk = ~clk;

wire  miss;
wire [31:0] rd_data;
reg  [31:0] index = 0, wr_data = 0, addr = 0;
reg  rd_req = 1'b0, wr_req = 1'b0;
reg rd_req_ff = 1'b0, miss_ff = 1'b0;
reg [31:0] validation_count = 0;

always @ (posedge clk or posedge rst)
    if(rst) begin
        rd_req_ff <= 1'b0;
        miss_ff   <= 1'b0;
    end else begin
        rd_req_ff <= rd_req;
        miss_ff   <= miss;
    end

always @ (posedge clk or posedge rst)
    if(rst) begin
        validation_count <= 0;
    end else begin
        if(validation_count>=`DATA_COUNT) begin
            validation_count <= 'hffffffff;
        end else if(rd_req_ff && (index>(4*`DATA_COUNT))) begin
            if(~miss_ff) begin
                if(validation_data[validation_count]==rd_data)
                    validation_count <= validation_count+1;
                else
                    validation_count <= 0;
            end
        end else begin
            validation_count <= 0;
        end
    end

always @ (posedge clk or posedge rst)
    if(rst) begin
        index   <= 0;
        wr_data <= 0;
        addr    <= 0;
        rd_req  <= 1'b0;
        wr_req  <= 1'b0;
    end else begin
        if(~miss) begin
            if(index<`RDWR_COUNT) begin
                if(wr_cycle[index]) begin
                    rd_req  <= 1'b0;
                    wr_req  <= 1'b1;
                end else if(rd_cycle[index]) begin
                    wr_data <= 0;
                    rd_req  <= 1'b1;
                    wr_req  <= 1'b0;
                end else begin
                    wr_data <= 0;
                    rd_req  <= 1'b0;
                    wr_req  <= 1'b0;
                end
                wr_data <= wr_data_rom[index];
                addr    <= addr_rom[index];
                index <= index + 1;
            end else begin
                wr_data <= 0;
                addr    <= 0;
                rd_req  <= 1'b0;
                wr_req  <= 1'b0;
            end
        end
    end

cache #(
    .LINE_ADDR_LEN  ( 3             ),
    .SET_ADDR_LEN   ( 2             ),
    .TAG_ADDR_LEN   ( 12            ),
    .WAY_CNT        ( 3             )
) cache_test_instance (
    .clk            ( clk           ),
    .rst            ( rst           ),
    .miss           ( miss          ),
    .addr           ( addr          ),
    .rd_req         ( rd_req        ),
    .rd_data        ( rd_data       ),
    .wr_req         ( wr_req        ),
    .wr_data        ( wr_data       )
);

endmodule

