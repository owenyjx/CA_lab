
module mem #(                   // 
    parameter  ADDR_LEN  = 11   // 
) (
    input  clk, rst,
    input  [ADDR_LEN-1:0] addr, // memory address
    output reg [31:0] rd_data,  // data read out
    input  wr_req,
    input  [31:0] wr_data       // data write in
);
localparam MEM_SIZE = 1<<ADDR_LEN;
reg [31:0] ram_cell [MEM_SIZE];

always @ (posedge clk or posedge rst)
    if(rst)
        rd_data <= 0;
    else
        rd_data <= ram_cell[addr];

always @ (posedge clk)
    if(wr_req) 
        ram_cell[addr] <= wr_data;

initial begin
    // dst matrix C
    ram_cell[       0] = 32'h0;  // 32'h20e1a6d5;
    ram_cell[       1] = 32'h0;  // 32'hf05e55d1;
    ram_cell[       2] = 32'h0;  // 32'h38b45bd7;
    ram_cell[       3] = 32'h0;  // 32'hc2eed978;
    ram_cell[       4] = 32'h0;  // 32'h8793e211;
    ram_cell[       5] = 32'h0;  // 32'h73bada01;
    ram_cell[       6] = 32'h0;  // 32'h676e0f68;
    ram_cell[       7] = 32'h0;  // 32'h2d0af092;
    ram_cell[       8] = 32'h0;  // 32'h066f22e5;
    ram_cell[       9] = 32'h0;  // 32'h7e2c4438;
    ram_cell[      10] = 32'h0;  // 32'h93c5a38a;
    ram_cell[      11] = 32'h0;  // 32'haf0fd0d5;
    ram_cell[      12] = 32'h0;  // 32'he422c3ac;
    ram_cell[      13] = 32'h0;  // 32'he88d7885;
    ram_cell[      14] = 32'h0;  // 32'h70c89105;
    ram_cell[      15] = 32'h0;  // 32'h94f06b22;
    ram_cell[      16] = 32'h0;  // 32'hd603257f;
    ram_cell[      17] = 32'h0;  // 32'h14452512;
    ram_cell[      18] = 32'h0;  // 32'h332a3c6e;
    ram_cell[      19] = 32'h0;  // 32'h16e4aa25;
    ram_cell[      20] = 32'h0;  // 32'h7e7df3ff;
    ram_cell[      21] = 32'h0;  // 32'h6de12f22;
    ram_cell[      22] = 32'h0;  // 32'h7b6ca402;
    ram_cell[      23] = 32'h0;  // 32'h355f1e55;
    ram_cell[      24] = 32'h0;  // 32'h8bde0bc9;
    ram_cell[      25] = 32'h0;  // 32'hcf98d45c;
    ram_cell[      26] = 32'h0;  // 32'h0fad9d88;
    ram_cell[      27] = 32'h0;  // 32'h443a5783;
    ram_cell[      28] = 32'h0;  // 32'hfa96d0ca;
    ram_cell[      29] = 32'h0;  // 32'h81c7ea22;
    ram_cell[      30] = 32'h0;  // 32'hcfdc0b3c;
    ram_cell[      31] = 32'h0;  // 32'hb045bc28;
    ram_cell[      32] = 32'h0;  // 32'h1c1985da;
    ram_cell[      33] = 32'h0;  // 32'hf38c9905;
    ram_cell[      34] = 32'h0;  // 32'h427e8d28;
    ram_cell[      35] = 32'h0;  // 32'hcd382712;
    ram_cell[      36] = 32'h0;  // 32'h476fea28;
    ram_cell[      37] = 32'h0;  // 32'hd7cfaf92;
    ram_cell[      38] = 32'h0;  // 32'h7cf66fd9;
    ram_cell[      39] = 32'h0;  // 32'h372192be;
    ram_cell[      40] = 32'h0;  // 32'h982a07b3;
    ram_cell[      41] = 32'h0;  // 32'hda1b72e5;
    ram_cell[      42] = 32'h0;  // 32'hb7bc972a;
    ram_cell[      43] = 32'h0;  // 32'h079284ec;
    ram_cell[      44] = 32'h0;  // 32'hadef499f;
    ram_cell[      45] = 32'h0;  // 32'h617b92d0;
    ram_cell[      46] = 32'h0;  // 32'h540d8a81;
    ram_cell[      47] = 32'h0;  // 32'had3ed61c;
    ram_cell[      48] = 32'h0;  // 32'hc8155869;
    ram_cell[      49] = 32'h0;  // 32'ha81e76b7;
    ram_cell[      50] = 32'h0;  // 32'h01adf758;
    ram_cell[      51] = 32'h0;  // 32'h13a9fe64;
    ram_cell[      52] = 32'h0;  // 32'h674e3c90;
    ram_cell[      53] = 32'h0;  // 32'h8c0482de;
    ram_cell[      54] = 32'h0;  // 32'h765b2d2f;
    ram_cell[      55] = 32'h0;  // 32'h0c3bd743;
    ram_cell[      56] = 32'h0;  // 32'he99c451e;
    ram_cell[      57] = 32'h0;  // 32'hb1048d88;
    ram_cell[      58] = 32'h0;  // 32'hec4c189d;
    ram_cell[      59] = 32'h0;  // 32'h06a5d237;
    ram_cell[      60] = 32'h0;  // 32'hb773c5fc;
    ram_cell[      61] = 32'h0;  // 32'haaeb03d0;
    ram_cell[      62] = 32'h0;  // 32'h5206a0e8;
    ram_cell[      63] = 32'h0;  // 32'hd3497b58;
    ram_cell[      64] = 32'h0;  // 32'h86801f9d;
    ram_cell[      65] = 32'h0;  // 32'h30e6a4c5;
    ram_cell[      66] = 32'h0;  // 32'h20782e2b;
    ram_cell[      67] = 32'h0;  // 32'hb92d8644;
    ram_cell[      68] = 32'h0;  // 32'h04477e03;
    ram_cell[      69] = 32'h0;  // 32'h95bec159;
    ram_cell[      70] = 32'h0;  // 32'h5250db52;
    ram_cell[      71] = 32'h0;  // 32'h79f94be5;
    ram_cell[      72] = 32'h0;  // 32'hd43f3955;
    ram_cell[      73] = 32'h0;  // 32'hde137ae6;
    ram_cell[      74] = 32'h0;  // 32'hbf1c785e;
    ram_cell[      75] = 32'h0;  // 32'h6ad14e66;
    ram_cell[      76] = 32'h0;  // 32'h63cc2d0b;
    ram_cell[      77] = 32'h0;  // 32'h28542acb;
    ram_cell[      78] = 32'h0;  // 32'h2befd856;
    ram_cell[      79] = 32'h0;  // 32'h790fb91b;
    ram_cell[      80] = 32'h0;  // 32'h65ff52b5;
    ram_cell[      81] = 32'h0;  // 32'hf2e9a9c2;
    ram_cell[      82] = 32'h0;  // 32'hf81d5510;
    ram_cell[      83] = 32'h0;  // 32'h62529759;
    ram_cell[      84] = 32'h0;  // 32'he743df09;
    ram_cell[      85] = 32'h0;  // 32'h8d53ec0b;
    ram_cell[      86] = 32'h0;  // 32'h753b8fb3;
    ram_cell[      87] = 32'h0;  // 32'hc26c4a0a;
    ram_cell[      88] = 32'h0;  // 32'h258e9dc4;
    ram_cell[      89] = 32'h0;  // 32'he23526f2;
    ram_cell[      90] = 32'h0;  // 32'h15308098;
    ram_cell[      91] = 32'h0;  // 32'h94c9a506;
    ram_cell[      92] = 32'h0;  // 32'h2452e8be;
    ram_cell[      93] = 32'h0;  // 32'hdaa592c6;
    ram_cell[      94] = 32'h0;  // 32'h8925a817;
    ram_cell[      95] = 32'h0;  // 32'hcee9e566;
    ram_cell[      96] = 32'h0;  // 32'hee891692;
    ram_cell[      97] = 32'h0;  // 32'hdf30e769;
    ram_cell[      98] = 32'h0;  // 32'h86f947fb;
    ram_cell[      99] = 32'h0;  // 32'h6a62eac1;
    ram_cell[     100] = 32'h0;  // 32'hb0a52b12;
    ram_cell[     101] = 32'h0;  // 32'h38f315e9;
    ram_cell[     102] = 32'h0;  // 32'h86cb0d4b;
    ram_cell[     103] = 32'h0;  // 32'hde83f933;
    ram_cell[     104] = 32'h0;  // 32'h6e0a906b;
    ram_cell[     105] = 32'h0;  // 32'ha45cdf31;
    ram_cell[     106] = 32'h0;  // 32'h27cbba85;
    ram_cell[     107] = 32'h0;  // 32'h2c418b08;
    ram_cell[     108] = 32'h0;  // 32'hb39e2936;
    ram_cell[     109] = 32'h0;  // 32'h7b4d938c;
    ram_cell[     110] = 32'h0;  // 32'h46b9d6f6;
    ram_cell[     111] = 32'h0;  // 32'h307da2f2;
    ram_cell[     112] = 32'h0;  // 32'hffbcb0d1;
    ram_cell[     113] = 32'h0;  // 32'h30aaa0e3;
    ram_cell[     114] = 32'h0;  // 32'h0cca938e;
    ram_cell[     115] = 32'h0;  // 32'hef7db367;
    ram_cell[     116] = 32'h0;  // 32'hf628450f;
    ram_cell[     117] = 32'h0;  // 32'h478654c1;
    ram_cell[     118] = 32'h0;  // 32'hf76888e4;
    ram_cell[     119] = 32'h0;  // 32'hc380629a;
    ram_cell[     120] = 32'h0;  // 32'h2ad48167;
    ram_cell[     121] = 32'h0;  // 32'h61d07951;
    ram_cell[     122] = 32'h0;  // 32'h8b35bf02;
    ram_cell[     123] = 32'h0;  // 32'hcd342b37;
    ram_cell[     124] = 32'h0;  // 32'hb1720e19;
    ram_cell[     125] = 32'h0;  // 32'h2bb26ce6;
    ram_cell[     126] = 32'h0;  // 32'hba58126e;
    ram_cell[     127] = 32'h0;  // 32'h9466a76e;
    ram_cell[     128] = 32'h0;  // 32'hc94a2dca;
    ram_cell[     129] = 32'h0;  // 32'h20c6052b;
    ram_cell[     130] = 32'h0;  // 32'h585fa1db;
    ram_cell[     131] = 32'h0;  // 32'he1d619d9;
    ram_cell[     132] = 32'h0;  // 32'h5c5937ed;
    ram_cell[     133] = 32'h0;  // 32'hb5ac42cd;
    ram_cell[     134] = 32'h0;  // 32'h311cd399;
    ram_cell[     135] = 32'h0;  // 32'hfd25a583;
    ram_cell[     136] = 32'h0;  // 32'h920d7e0c;
    ram_cell[     137] = 32'h0;  // 32'h8a5fd4c8;
    ram_cell[     138] = 32'h0;  // 32'h8093de5d;
    ram_cell[     139] = 32'h0;  // 32'h6fc123e7;
    ram_cell[     140] = 32'h0;  // 32'hb7f2492d;
    ram_cell[     141] = 32'h0;  // 32'hea9640ad;
    ram_cell[     142] = 32'h0;  // 32'h36057091;
    ram_cell[     143] = 32'h0;  // 32'h11c92065;
    ram_cell[     144] = 32'h0;  // 32'h0460005d;
    ram_cell[     145] = 32'h0;  // 32'h21817731;
    ram_cell[     146] = 32'h0;  // 32'h0294043c;
    ram_cell[     147] = 32'h0;  // 32'h0acbf7eb;
    ram_cell[     148] = 32'h0;  // 32'h185e2e75;
    ram_cell[     149] = 32'h0;  // 32'ha31e9a62;
    ram_cell[     150] = 32'h0;  // 32'h51afd841;
    ram_cell[     151] = 32'h0;  // 32'h0c27bd45;
    ram_cell[     152] = 32'h0;  // 32'h48ce773e;
    ram_cell[     153] = 32'h0;  // 32'h70bc982a;
    ram_cell[     154] = 32'h0;  // 32'h44088baa;
    ram_cell[     155] = 32'h0;  // 32'hbcd53900;
    ram_cell[     156] = 32'h0;  // 32'hbd07a9c2;
    ram_cell[     157] = 32'h0;  // 32'h10f7c950;
    ram_cell[     158] = 32'h0;  // 32'hc60607ae;
    ram_cell[     159] = 32'h0;  // 32'hadd11700;
    ram_cell[     160] = 32'h0;  // 32'h4d922202;
    ram_cell[     161] = 32'h0;  // 32'hac619d8c;
    ram_cell[     162] = 32'h0;  // 32'hc0893b07;
    ram_cell[     163] = 32'h0;  // 32'h1982e763;
    ram_cell[     164] = 32'h0;  // 32'h05231243;
    ram_cell[     165] = 32'h0;  // 32'h76013682;
    ram_cell[     166] = 32'h0;  // 32'h52ab94f3;
    ram_cell[     167] = 32'h0;  // 32'h224989f2;
    ram_cell[     168] = 32'h0;  // 32'hc1a8a443;
    ram_cell[     169] = 32'h0;  // 32'h1eb1a5d4;
    ram_cell[     170] = 32'h0;  // 32'ha69e173a;
    ram_cell[     171] = 32'h0;  // 32'h792ecf58;
    ram_cell[     172] = 32'h0;  // 32'h452b01cc;
    ram_cell[     173] = 32'h0;  // 32'h870df736;
    ram_cell[     174] = 32'h0;  // 32'h14e522a6;
    ram_cell[     175] = 32'h0;  // 32'h87103aec;
    ram_cell[     176] = 32'h0;  // 32'h6d7cd5e1;
    ram_cell[     177] = 32'h0;  // 32'he6bd39f8;
    ram_cell[     178] = 32'h0;  // 32'h7c9e0af2;
    ram_cell[     179] = 32'h0;  // 32'hcb3cfcbb;
    ram_cell[     180] = 32'h0;  // 32'h0d6048e2;
    ram_cell[     181] = 32'h0;  // 32'hcf6a9abd;
    ram_cell[     182] = 32'h0;  // 32'h0a5637e7;
    ram_cell[     183] = 32'h0;  // 32'hb9b31346;
    ram_cell[     184] = 32'h0;  // 32'hae376a50;
    ram_cell[     185] = 32'h0;  // 32'hc3346e75;
    ram_cell[     186] = 32'h0;  // 32'ha4badbe8;
    ram_cell[     187] = 32'h0;  // 32'h0102426c;
    ram_cell[     188] = 32'h0;  // 32'ha61330f5;
    ram_cell[     189] = 32'h0;  // 32'hfcbc56c3;
    ram_cell[     190] = 32'h0;  // 32'h087600df;
    ram_cell[     191] = 32'h0;  // 32'hf4c2b90e;
    ram_cell[     192] = 32'h0;  // 32'hcb627241;
    ram_cell[     193] = 32'h0;  // 32'hb9dc354e;
    ram_cell[     194] = 32'h0;  // 32'hfd41ab03;
    ram_cell[     195] = 32'h0;  // 32'h895b9b46;
    ram_cell[     196] = 32'h0;  // 32'h365e08ec;
    ram_cell[     197] = 32'h0;  // 32'hd7bdfc5d;
    ram_cell[     198] = 32'h0;  // 32'he7e94735;
    ram_cell[     199] = 32'h0;  // 32'h13ee746f;
    ram_cell[     200] = 32'h0;  // 32'h73a50726;
    ram_cell[     201] = 32'h0;  // 32'ha6d50a27;
    ram_cell[     202] = 32'h0;  // 32'ha0bfd246;
    ram_cell[     203] = 32'h0;  // 32'ha9dfa92d;
    ram_cell[     204] = 32'h0;  // 32'h00a97e04;
    ram_cell[     205] = 32'h0;  // 32'h84b006bf;
    ram_cell[     206] = 32'h0;  // 32'h69bb3174;
    ram_cell[     207] = 32'h0;  // 32'hc20a3f60;
    ram_cell[     208] = 32'h0;  // 32'hb58e4496;
    ram_cell[     209] = 32'h0;  // 32'h5931ddf9;
    ram_cell[     210] = 32'h0;  // 32'h51c2d37b;
    ram_cell[     211] = 32'h0;  // 32'h26a0e22e;
    ram_cell[     212] = 32'h0;  // 32'h2ec42bdc;
    ram_cell[     213] = 32'h0;  // 32'h805e560e;
    ram_cell[     214] = 32'h0;  // 32'h49aead93;
    ram_cell[     215] = 32'h0;  // 32'hf2c07353;
    ram_cell[     216] = 32'h0;  // 32'hda846b52;
    ram_cell[     217] = 32'h0;  // 32'h80d380c5;
    ram_cell[     218] = 32'h0;  // 32'he0f46ba6;
    ram_cell[     219] = 32'h0;  // 32'hd43cf91b;
    ram_cell[     220] = 32'h0;  // 32'hcd5961b4;
    ram_cell[     221] = 32'h0;  // 32'h8cc84375;
    ram_cell[     222] = 32'h0;  // 32'haff5d9e1;
    ram_cell[     223] = 32'h0;  // 32'h82b91ca3;
    ram_cell[     224] = 32'h0;  // 32'h1c297b45;
    ram_cell[     225] = 32'h0;  // 32'h0826a9b6;
    ram_cell[     226] = 32'h0;  // 32'h6020fe6f;
    ram_cell[     227] = 32'h0;  // 32'he18e0ef9;
    ram_cell[     228] = 32'h0;  // 32'ha0295e49;
    ram_cell[     229] = 32'h0;  // 32'h773eefda;
    ram_cell[     230] = 32'h0;  // 32'ha900ea75;
    ram_cell[     231] = 32'h0;  // 32'h5391951d;
    ram_cell[     232] = 32'h0;  // 32'h78d57325;
    ram_cell[     233] = 32'h0;  // 32'h97729712;
    ram_cell[     234] = 32'h0;  // 32'h746e3f30;
    ram_cell[     235] = 32'h0;  // 32'h1f787187;
    ram_cell[     236] = 32'h0;  // 32'h328f44c6;
    ram_cell[     237] = 32'h0;  // 32'h09f21a27;
    ram_cell[     238] = 32'h0;  // 32'h38fc729e;
    ram_cell[     239] = 32'h0;  // 32'hbda53d37;
    ram_cell[     240] = 32'h0;  // 32'h6ed1b6a4;
    ram_cell[     241] = 32'h0;  // 32'hbfb8821a;
    ram_cell[     242] = 32'h0;  // 32'h4c97241f;
    ram_cell[     243] = 32'h0;  // 32'hdb608f2e;
    ram_cell[     244] = 32'h0;  // 32'ha3c98290;
    ram_cell[     245] = 32'h0;  // 32'h970765a0;
    ram_cell[     246] = 32'h0;  // 32'h73d8d704;
    ram_cell[     247] = 32'h0;  // 32'ha18325fc;
    ram_cell[     248] = 32'h0;  // 32'h71065bc2;
    ram_cell[     249] = 32'h0;  // 32'hcf8c751f;
    ram_cell[     250] = 32'h0;  // 32'hd9409775;
    ram_cell[     251] = 32'h0;  // 32'h699fb1bd;
    ram_cell[     252] = 32'h0;  // 32'h1707383e;
    ram_cell[     253] = 32'h0;  // 32'h152885a6;
    ram_cell[     254] = 32'h0;  // 32'hdbd3330c;
    ram_cell[     255] = 32'h0;  // 32'h3c2452b9;
    // src matrix A
    ram_cell[     256] = 32'h8e8731ff;
    ram_cell[     257] = 32'h06f3ffcf;
    ram_cell[     258] = 32'h8a9aeb42;
    ram_cell[     259] = 32'h21251d8f;
    ram_cell[     260] = 32'hc3ee7e9a;
    ram_cell[     261] = 32'h6244f464;
    ram_cell[     262] = 32'h8a871a23;
    ram_cell[     263] = 32'h52f72c54;
    ram_cell[     264] = 32'h0efc2dd6;
    ram_cell[     265] = 32'hb8a5a972;
    ram_cell[     266] = 32'h6d78a9d9;
    ram_cell[     267] = 32'hfb1144e6;
    ram_cell[     268] = 32'h1481a672;
    ram_cell[     269] = 32'h2a4230b0;
    ram_cell[     270] = 32'hab383dbc;
    ram_cell[     271] = 32'h18c5e7eb;
    ram_cell[     272] = 32'h33c5d12c;
    ram_cell[     273] = 32'h5a0c1cc0;
    ram_cell[     274] = 32'h41c91ff7;
    ram_cell[     275] = 32'h397b2e72;
    ram_cell[     276] = 32'h9113f90c;
    ram_cell[     277] = 32'h96840bc2;
    ram_cell[     278] = 32'h8e72eaca;
    ram_cell[     279] = 32'h61ba9053;
    ram_cell[     280] = 32'h2b064455;
    ram_cell[     281] = 32'h0f143e80;
    ram_cell[     282] = 32'hf0454641;
    ram_cell[     283] = 32'h6f94a4a3;
    ram_cell[     284] = 32'hb0f4e66c;
    ram_cell[     285] = 32'hd3fbfacb;
    ram_cell[     286] = 32'h825c21bb;
    ram_cell[     287] = 32'h605448d4;
    ram_cell[     288] = 32'h35c1bc0b;
    ram_cell[     289] = 32'hcd8fd09f;
    ram_cell[     290] = 32'hc57898ff;
    ram_cell[     291] = 32'hba2174f1;
    ram_cell[     292] = 32'h14270bbe;
    ram_cell[     293] = 32'h692f103f;
    ram_cell[     294] = 32'hce7039bf;
    ram_cell[     295] = 32'h68114852;
    ram_cell[     296] = 32'h00e8eb07;
    ram_cell[     297] = 32'ha8711320;
    ram_cell[     298] = 32'h0a8ee9ba;
    ram_cell[     299] = 32'hb44a4c7c;
    ram_cell[     300] = 32'hd10f0b6a;
    ram_cell[     301] = 32'hc3a13149;
    ram_cell[     302] = 32'h6c725dd5;
    ram_cell[     303] = 32'hddfe0a34;
    ram_cell[     304] = 32'h09890fb6;
    ram_cell[     305] = 32'hd08a18b2;
    ram_cell[     306] = 32'hc4e8960f;
    ram_cell[     307] = 32'he4f8aaf5;
    ram_cell[     308] = 32'h24b46316;
    ram_cell[     309] = 32'hd56dac8e;
    ram_cell[     310] = 32'h02f185d9;
    ram_cell[     311] = 32'h3e24dea9;
    ram_cell[     312] = 32'h2b443da3;
    ram_cell[     313] = 32'he374e4dc;
    ram_cell[     314] = 32'he2138055;
    ram_cell[     315] = 32'h1ee155a7;
    ram_cell[     316] = 32'h25c98e07;
    ram_cell[     317] = 32'hef9e60d9;
    ram_cell[     318] = 32'h320db41f;
    ram_cell[     319] = 32'h180f44d5;
    ram_cell[     320] = 32'h743a9004;
    ram_cell[     321] = 32'h11ae25d4;
    ram_cell[     322] = 32'h1e45daf7;
    ram_cell[     323] = 32'h56e63839;
    ram_cell[     324] = 32'h31bec569;
    ram_cell[     325] = 32'h28c7ba3a;
    ram_cell[     326] = 32'h32dce278;
    ram_cell[     327] = 32'h1f59f793;
    ram_cell[     328] = 32'h979edd2d;
    ram_cell[     329] = 32'h2019b7ca;
    ram_cell[     330] = 32'h1f18f78d;
    ram_cell[     331] = 32'hbfdc1768;
    ram_cell[     332] = 32'hc6b5ff69;
    ram_cell[     333] = 32'h7c8b0e3d;
    ram_cell[     334] = 32'h28aaf320;
    ram_cell[     335] = 32'h6dc37373;
    ram_cell[     336] = 32'h4517b609;
    ram_cell[     337] = 32'h32438e59;
    ram_cell[     338] = 32'h6ad4cf3c;
    ram_cell[     339] = 32'h0218310b;
    ram_cell[     340] = 32'hfe857164;
    ram_cell[     341] = 32'hd982b5a6;
    ram_cell[     342] = 32'h63aeabb9;
    ram_cell[     343] = 32'hca72b858;
    ram_cell[     344] = 32'h5b2ff645;
    ram_cell[     345] = 32'ha270b32b;
    ram_cell[     346] = 32'h8bef048c;
    ram_cell[     347] = 32'h1ad43d47;
    ram_cell[     348] = 32'hc8a72ccb;
    ram_cell[     349] = 32'hb5203436;
    ram_cell[     350] = 32'h61302cc2;
    ram_cell[     351] = 32'h1c5f1619;
    ram_cell[     352] = 32'h47e60e0e;
    ram_cell[     353] = 32'hefcd79e7;
    ram_cell[     354] = 32'hd1136752;
    ram_cell[     355] = 32'h3813441b;
    ram_cell[     356] = 32'ha2ff648c;
    ram_cell[     357] = 32'h5851f387;
    ram_cell[     358] = 32'hdc6f0100;
    ram_cell[     359] = 32'h53526ce2;
    ram_cell[     360] = 32'h81be7902;
    ram_cell[     361] = 32'hc01e42cb;
    ram_cell[     362] = 32'he79f40e6;
    ram_cell[     363] = 32'h6a35d3df;
    ram_cell[     364] = 32'he47daf9b;
    ram_cell[     365] = 32'hc36dacf2;
    ram_cell[     366] = 32'he66eae50;
    ram_cell[     367] = 32'h98c4b046;
    ram_cell[     368] = 32'h1da2b65a;
    ram_cell[     369] = 32'h2b2f8783;
    ram_cell[     370] = 32'hebafd47a;
    ram_cell[     371] = 32'ha07fa5dd;
    ram_cell[     372] = 32'hfe648b31;
    ram_cell[     373] = 32'h6815e14f;
    ram_cell[     374] = 32'hf87b5bf6;
    ram_cell[     375] = 32'h87ec21c9;
    ram_cell[     376] = 32'h9f2bad7a;
    ram_cell[     377] = 32'hecd9d7f8;
    ram_cell[     378] = 32'h8f995e4f;
    ram_cell[     379] = 32'hdb812200;
    ram_cell[     380] = 32'h734c872e;
    ram_cell[     381] = 32'hd5880abd;
    ram_cell[     382] = 32'hcd80a051;
    ram_cell[     383] = 32'h35eeb5f0;
    ram_cell[     384] = 32'hf7011394;
    ram_cell[     385] = 32'hc20ddb67;
    ram_cell[     386] = 32'h784a4e18;
    ram_cell[     387] = 32'hf6817f85;
    ram_cell[     388] = 32'h30a31e3f;
    ram_cell[     389] = 32'h2f9f8b88;
    ram_cell[     390] = 32'hdbc9b96a;
    ram_cell[     391] = 32'h4e1c536e;
    ram_cell[     392] = 32'h8cd16562;
    ram_cell[     393] = 32'hbdff36b8;
    ram_cell[     394] = 32'hbd56512a;
    ram_cell[     395] = 32'he147f66f;
    ram_cell[     396] = 32'hdcf353c3;
    ram_cell[     397] = 32'hf9ef7965;
    ram_cell[     398] = 32'hc17cf791;
    ram_cell[     399] = 32'hd4299ed0;
    ram_cell[     400] = 32'h65b8bcbe;
    ram_cell[     401] = 32'h2fbc6d09;
    ram_cell[     402] = 32'h1ffb8266;
    ram_cell[     403] = 32'h2125699a;
    ram_cell[     404] = 32'hae4ee5a2;
    ram_cell[     405] = 32'h0f36e496;
    ram_cell[     406] = 32'h3225123c;
    ram_cell[     407] = 32'h8069c91d;
    ram_cell[     408] = 32'ha174d88e;
    ram_cell[     409] = 32'hc943130d;
    ram_cell[     410] = 32'h9b0ddd20;
    ram_cell[     411] = 32'hfd57f195;
    ram_cell[     412] = 32'h9101a45a;
    ram_cell[     413] = 32'h49428f8a;
    ram_cell[     414] = 32'h9462fe80;
    ram_cell[     415] = 32'h81831b50;
    ram_cell[     416] = 32'he732c135;
    ram_cell[     417] = 32'h12463b77;
    ram_cell[     418] = 32'h27634c25;
    ram_cell[     419] = 32'h3c84d9c9;
    ram_cell[     420] = 32'h16e74561;
    ram_cell[     421] = 32'h0d22356e;
    ram_cell[     422] = 32'he52feab7;
    ram_cell[     423] = 32'h22c36f72;
    ram_cell[     424] = 32'h9a75d836;
    ram_cell[     425] = 32'h0097ba5d;
    ram_cell[     426] = 32'hd2dacdcf;
    ram_cell[     427] = 32'hd03aac55;
    ram_cell[     428] = 32'h06fe61c9;
    ram_cell[     429] = 32'h5f517737;
    ram_cell[     430] = 32'hc20c3b8c;
    ram_cell[     431] = 32'h0cc94165;
    ram_cell[     432] = 32'hc7960a7c;
    ram_cell[     433] = 32'h413c34b8;
    ram_cell[     434] = 32'h1e48b581;
    ram_cell[     435] = 32'h76f8c8d9;
    ram_cell[     436] = 32'h918c8207;
    ram_cell[     437] = 32'h110fa994;
    ram_cell[     438] = 32'h7d6b01ee;
    ram_cell[     439] = 32'h7173a186;
    ram_cell[     440] = 32'h4cba53a0;
    ram_cell[     441] = 32'haacd1388;
    ram_cell[     442] = 32'he65c59a4;
    ram_cell[     443] = 32'h2a66b087;
    ram_cell[     444] = 32'h2072e249;
    ram_cell[     445] = 32'hc39c865c;
    ram_cell[     446] = 32'h14db6c45;
    ram_cell[     447] = 32'ha816f161;
    ram_cell[     448] = 32'h0611d9c5;
    ram_cell[     449] = 32'h133969e9;
    ram_cell[     450] = 32'he6dcbb05;
    ram_cell[     451] = 32'h6ae11072;
    ram_cell[     452] = 32'hc009f409;
    ram_cell[     453] = 32'hfd8cbd73;
    ram_cell[     454] = 32'h11ac73ba;
    ram_cell[     455] = 32'h0f673680;
    ram_cell[     456] = 32'h69405a0d;
    ram_cell[     457] = 32'h9634e5d3;
    ram_cell[     458] = 32'h34cccc8c;
    ram_cell[     459] = 32'h8ffef50d;
    ram_cell[     460] = 32'h0cc15efc;
    ram_cell[     461] = 32'h71b1db4d;
    ram_cell[     462] = 32'hac053979;
    ram_cell[     463] = 32'ha3abf277;
    ram_cell[     464] = 32'hc73244ea;
    ram_cell[     465] = 32'h1397b4bc;
    ram_cell[     466] = 32'h6d7c4818;
    ram_cell[     467] = 32'hc3fb78e4;
    ram_cell[     468] = 32'h38da019f;
    ram_cell[     469] = 32'h1bbef8de;
    ram_cell[     470] = 32'haf696594;
    ram_cell[     471] = 32'h75e58fc0;
    ram_cell[     472] = 32'hba6f81c0;
    ram_cell[     473] = 32'hcf170095;
    ram_cell[     474] = 32'h71bb1920;
    ram_cell[     475] = 32'h5287418b;
    ram_cell[     476] = 32'hbcb75b41;
    ram_cell[     477] = 32'h7526bdd3;
    ram_cell[     478] = 32'heb71e905;
    ram_cell[     479] = 32'h2cc92b1b;
    ram_cell[     480] = 32'hd1978fc0;
    ram_cell[     481] = 32'h30e5a950;
    ram_cell[     482] = 32'h4effd79f;
    ram_cell[     483] = 32'hf18fe14a;
    ram_cell[     484] = 32'h6849fe29;
    ram_cell[     485] = 32'h0b315010;
    ram_cell[     486] = 32'hbea3e15c;
    ram_cell[     487] = 32'ha34f7911;
    ram_cell[     488] = 32'h642ba777;
    ram_cell[     489] = 32'hf6b6829a;
    ram_cell[     490] = 32'h3f402424;
    ram_cell[     491] = 32'h9c5049d3;
    ram_cell[     492] = 32'ha31100ba;
    ram_cell[     493] = 32'h560d2115;
    ram_cell[     494] = 32'h4f0b3191;
    ram_cell[     495] = 32'hfe61e1e5;
    ram_cell[     496] = 32'hb8d1deab;
    ram_cell[     497] = 32'h100474e1;
    ram_cell[     498] = 32'h08d5e81e;
    ram_cell[     499] = 32'he4ae6620;
    ram_cell[     500] = 32'hb1f1289d;
    ram_cell[     501] = 32'h7d47259c;
    ram_cell[     502] = 32'hfc383a23;
    ram_cell[     503] = 32'h82bf3617;
    ram_cell[     504] = 32'h5cb516a9;
    ram_cell[     505] = 32'h9410c732;
    ram_cell[     506] = 32'h83ca3b53;
    ram_cell[     507] = 32'hcb674f7e;
    ram_cell[     508] = 32'hf1856362;
    ram_cell[     509] = 32'hdffc5b7b;
    ram_cell[     510] = 32'h6aae8e61;
    ram_cell[     511] = 32'h926e9862;
    // src matrix B
    ram_cell[     512] = 32'h6f8a6e0d;
    ram_cell[     513] = 32'h2464b7ae;
    ram_cell[     514] = 32'h7550e19f;
    ram_cell[     515] = 32'h37293236;
    ram_cell[     516] = 32'h4ad6dfba;
    ram_cell[     517] = 32'hee33d05c;
    ram_cell[     518] = 32'h3483d1a5;
    ram_cell[     519] = 32'h4ea13038;
    ram_cell[     520] = 32'h7371e24a;
    ram_cell[     521] = 32'hfa84eb1f;
    ram_cell[     522] = 32'h51065496;
    ram_cell[     523] = 32'h889f3d6c;
    ram_cell[     524] = 32'hceafcf7e;
    ram_cell[     525] = 32'hb3e7869b;
    ram_cell[     526] = 32'hd9ac4196;
    ram_cell[     527] = 32'h01f8acb2;
    ram_cell[     528] = 32'h5deeaa5f;
    ram_cell[     529] = 32'h784b71d2;
    ram_cell[     530] = 32'h520e9363;
    ram_cell[     531] = 32'h53f621b0;
    ram_cell[     532] = 32'h4537453d;
    ram_cell[     533] = 32'h954ef7ad;
    ram_cell[     534] = 32'hfe9498a5;
    ram_cell[     535] = 32'h2f07fbf1;
    ram_cell[     536] = 32'ha795744d;
    ram_cell[     537] = 32'hddb88b62;
    ram_cell[     538] = 32'h2a497871;
    ram_cell[     539] = 32'ha4bd4128;
    ram_cell[     540] = 32'hb5d96d58;
    ram_cell[     541] = 32'h74f30a68;
    ram_cell[     542] = 32'h7a0dd32b;
    ram_cell[     543] = 32'h1dc4deff;
    ram_cell[     544] = 32'hfbdb71dd;
    ram_cell[     545] = 32'h6aa06b2d;
    ram_cell[     546] = 32'h71f2fcdf;
    ram_cell[     547] = 32'hc1002f28;
    ram_cell[     548] = 32'hf12fc996;
    ram_cell[     549] = 32'hb10a960e;
    ram_cell[     550] = 32'h04010845;
    ram_cell[     551] = 32'h9c8f898a;
    ram_cell[     552] = 32'h501ef374;
    ram_cell[     553] = 32'hd855e433;
    ram_cell[     554] = 32'hfbc1948a;
    ram_cell[     555] = 32'hcf84af1b;
    ram_cell[     556] = 32'h5a0db9b8;
    ram_cell[     557] = 32'h146bdaa6;
    ram_cell[     558] = 32'he48d79b5;
    ram_cell[     559] = 32'h75cd0027;
    ram_cell[     560] = 32'h61f5eea0;
    ram_cell[     561] = 32'h0e9f8b6e;
    ram_cell[     562] = 32'hb8bbb359;
    ram_cell[     563] = 32'h55081b47;
    ram_cell[     564] = 32'hdf620bff;
    ram_cell[     565] = 32'he7d32cee;
    ram_cell[     566] = 32'h96a229c9;
    ram_cell[     567] = 32'hfb6d6f72;
    ram_cell[     568] = 32'hd083306b;
    ram_cell[     569] = 32'hecfe65e8;
    ram_cell[     570] = 32'h7b78bd25;
    ram_cell[     571] = 32'h0c7ef6e3;
    ram_cell[     572] = 32'h7989b850;
    ram_cell[     573] = 32'ha2cfa710;
    ram_cell[     574] = 32'haddf1ac6;
    ram_cell[     575] = 32'h52abc981;
    ram_cell[     576] = 32'hebc23bdb;
    ram_cell[     577] = 32'hba654a0c;
    ram_cell[     578] = 32'h82b6551a;
    ram_cell[     579] = 32'hc8b47ba1;
    ram_cell[     580] = 32'h678ec5fa;
    ram_cell[     581] = 32'h0be08731;
    ram_cell[     582] = 32'h498b2e15;
    ram_cell[     583] = 32'h45909f87;
    ram_cell[     584] = 32'h453228f3;
    ram_cell[     585] = 32'h46b34275;
    ram_cell[     586] = 32'h0eb53a5a;
    ram_cell[     587] = 32'hebd48305;
    ram_cell[     588] = 32'h1cc02db9;
    ram_cell[     589] = 32'had3c1278;
    ram_cell[     590] = 32'h68ae12e2;
    ram_cell[     591] = 32'h86f6a419;
    ram_cell[     592] = 32'h11717f2b;
    ram_cell[     593] = 32'h80fb7081;
    ram_cell[     594] = 32'h38599c8a;
    ram_cell[     595] = 32'hfaf1dbbe;
    ram_cell[     596] = 32'h79ea385b;
    ram_cell[     597] = 32'h9646e4b4;
    ram_cell[     598] = 32'hbad69c39;
    ram_cell[     599] = 32'h1d46cc82;
    ram_cell[     600] = 32'hc34bb886;
    ram_cell[     601] = 32'h2dde108e;
    ram_cell[     602] = 32'hf368a724;
    ram_cell[     603] = 32'he15b4a55;
    ram_cell[     604] = 32'h008b4432;
    ram_cell[     605] = 32'he0f742bd;
    ram_cell[     606] = 32'h98d2ef26;
    ram_cell[     607] = 32'h7c774d7d;
    ram_cell[     608] = 32'h8fc50efe;
    ram_cell[     609] = 32'h9785544b;
    ram_cell[     610] = 32'h1ba82293;
    ram_cell[     611] = 32'hc38b5b4c;
    ram_cell[     612] = 32'h4bee192d;
    ram_cell[     613] = 32'hae93ef95;
    ram_cell[     614] = 32'h97215021;
    ram_cell[     615] = 32'h5560f4da;
    ram_cell[     616] = 32'hd06f06ca;
    ram_cell[     617] = 32'h72817b1c;
    ram_cell[     618] = 32'h12eb41ec;
    ram_cell[     619] = 32'h5754e0e1;
    ram_cell[     620] = 32'hae43f57b;
    ram_cell[     621] = 32'ha3d3a7b3;
    ram_cell[     622] = 32'h7c9d9e50;
    ram_cell[     623] = 32'h6d785bde;
    ram_cell[     624] = 32'ha05f04be;
    ram_cell[     625] = 32'h0ff4e385;
    ram_cell[     626] = 32'h90497dff;
    ram_cell[     627] = 32'h6789706f;
    ram_cell[     628] = 32'h8ec254f9;
    ram_cell[     629] = 32'hc9d8824b;
    ram_cell[     630] = 32'h368a0f0c;
    ram_cell[     631] = 32'hdd067e3d;
    ram_cell[     632] = 32'h95e9ced5;
    ram_cell[     633] = 32'h1c20c9d2;
    ram_cell[     634] = 32'h029405c1;
    ram_cell[     635] = 32'h4a4ff995;
    ram_cell[     636] = 32'h82de4966;
    ram_cell[     637] = 32'h305c94e4;
    ram_cell[     638] = 32'h38665993;
    ram_cell[     639] = 32'h1a92cca3;
    ram_cell[     640] = 32'h3b6afc5b;
    ram_cell[     641] = 32'h03f92849;
    ram_cell[     642] = 32'h80269072;
    ram_cell[     643] = 32'h6bd2c23e;
    ram_cell[     644] = 32'hbece464c;
    ram_cell[     645] = 32'h745924d4;
    ram_cell[     646] = 32'h3bbc1a08;
    ram_cell[     647] = 32'h4d25c556;
    ram_cell[     648] = 32'h53d9c88a;
    ram_cell[     649] = 32'h871eea93;
    ram_cell[     650] = 32'hf9c954ae;
    ram_cell[     651] = 32'h2d89ccf7;
    ram_cell[     652] = 32'h4a128004;
    ram_cell[     653] = 32'h863dde97;
    ram_cell[     654] = 32'h471b9e26;
    ram_cell[     655] = 32'hd55f8a17;
    ram_cell[     656] = 32'h269099ad;
    ram_cell[     657] = 32'h927d7b66;
    ram_cell[     658] = 32'h6bb605e5;
    ram_cell[     659] = 32'hf830baea;
    ram_cell[     660] = 32'h3792196e;
    ram_cell[     661] = 32'hfca4fb93;
    ram_cell[     662] = 32'h947b2ddb;
    ram_cell[     663] = 32'h229435b0;
    ram_cell[     664] = 32'h9cb8373f;
    ram_cell[     665] = 32'hc242bd48;
    ram_cell[     666] = 32'hd55c1dfc;
    ram_cell[     667] = 32'hdab97dce;
    ram_cell[     668] = 32'h27e7f6bc;
    ram_cell[     669] = 32'h814b8d5e;
    ram_cell[     670] = 32'hb7d3a0a6;
    ram_cell[     671] = 32'h0d956ec8;
    ram_cell[     672] = 32'h5dbfa9a3;
    ram_cell[     673] = 32'hbe212e24;
    ram_cell[     674] = 32'h445d37be;
    ram_cell[     675] = 32'h8a0639d7;
    ram_cell[     676] = 32'hde57e4fd;
    ram_cell[     677] = 32'hfab08850;
    ram_cell[     678] = 32'hdfc696a7;
    ram_cell[     679] = 32'h992d40a6;
    ram_cell[     680] = 32'ha9f1c8d2;
    ram_cell[     681] = 32'h9c501c32;
    ram_cell[     682] = 32'h2f0fb23d;
    ram_cell[     683] = 32'hac9d32b8;
    ram_cell[     684] = 32'hcacb062c;
    ram_cell[     685] = 32'h541cfff5;
    ram_cell[     686] = 32'ha15422a7;
    ram_cell[     687] = 32'h7d2dd3a6;
    ram_cell[     688] = 32'h53b3c5dd;
    ram_cell[     689] = 32'hf18a4f08;
    ram_cell[     690] = 32'hbbc6e4c7;
    ram_cell[     691] = 32'h44f777e6;
    ram_cell[     692] = 32'h80664f6d;
    ram_cell[     693] = 32'h9350580d;
    ram_cell[     694] = 32'h0230f03b;
    ram_cell[     695] = 32'h8490b933;
    ram_cell[     696] = 32'h5e263b03;
    ram_cell[     697] = 32'h1c3eeb56;
    ram_cell[     698] = 32'h7345e8c2;
    ram_cell[     699] = 32'h6d444f2b;
    ram_cell[     700] = 32'h9c9a0b46;
    ram_cell[     701] = 32'h73ab1cac;
    ram_cell[     702] = 32'h404b0fcc;
    ram_cell[     703] = 32'h20c4d3e2;
    ram_cell[     704] = 32'h878edcb6;
    ram_cell[     705] = 32'h8f5e5716;
    ram_cell[     706] = 32'h0351c7f5;
    ram_cell[     707] = 32'h551dced6;
    ram_cell[     708] = 32'h432be16e;
    ram_cell[     709] = 32'h044d2ab0;
    ram_cell[     710] = 32'h1e1dcc40;
    ram_cell[     711] = 32'h4fffe765;
    ram_cell[     712] = 32'h12ea7ee9;
    ram_cell[     713] = 32'h870476b7;
    ram_cell[     714] = 32'hf12bf54f;
    ram_cell[     715] = 32'h1542aca3;
    ram_cell[     716] = 32'h66b0eabc;
    ram_cell[     717] = 32'h04724ef5;
    ram_cell[     718] = 32'h8a7c12fd;
    ram_cell[     719] = 32'h1d97b181;
    ram_cell[     720] = 32'h386b409b;
    ram_cell[     721] = 32'h021998fe;
    ram_cell[     722] = 32'hea1720e6;
    ram_cell[     723] = 32'h0574da7c;
    ram_cell[     724] = 32'hc0fa7e83;
    ram_cell[     725] = 32'hd4df5372;
    ram_cell[     726] = 32'hbe7c4373;
    ram_cell[     727] = 32'h9b74cf4d;
    ram_cell[     728] = 32'h391dee6c;
    ram_cell[     729] = 32'h99dce885;
    ram_cell[     730] = 32'h8f19515b;
    ram_cell[     731] = 32'he99c8dcb;
    ram_cell[     732] = 32'h54a93113;
    ram_cell[     733] = 32'hc025964a;
    ram_cell[     734] = 32'h3488aeeb;
    ram_cell[     735] = 32'h37db0c11;
    ram_cell[     736] = 32'h12aaea52;
    ram_cell[     737] = 32'h6335df39;
    ram_cell[     738] = 32'h42f28713;
    ram_cell[     739] = 32'h2948ac3b;
    ram_cell[     740] = 32'h3a797f43;
    ram_cell[     741] = 32'he2f4e670;
    ram_cell[     742] = 32'h6bfd1e5a;
    ram_cell[     743] = 32'h10aea374;
    ram_cell[     744] = 32'h928cb4cb;
    ram_cell[     745] = 32'h463f5e65;
    ram_cell[     746] = 32'h298f1623;
    ram_cell[     747] = 32'hb860f2ee;
    ram_cell[     748] = 32'hc8d9f347;
    ram_cell[     749] = 32'h8f236a32;
    ram_cell[     750] = 32'hbab04c60;
    ram_cell[     751] = 32'he8bd1fd0;
    ram_cell[     752] = 32'h7dc37944;
    ram_cell[     753] = 32'ha21d72a8;
    ram_cell[     754] = 32'he53b9b19;
    ram_cell[     755] = 32'hcbc5f4fe;
    ram_cell[     756] = 32'h13922ebd;
    ram_cell[     757] = 32'hd3487a4d;
    ram_cell[     758] = 32'h936af2b7;
    ram_cell[     759] = 32'hff7b2145;
    ram_cell[     760] = 32'h75348e99;
    ram_cell[     761] = 32'h3b67c8ef;
    ram_cell[     762] = 32'h0421f3db;
    ram_cell[     763] = 32'h379ac443;
    ram_cell[     764] = 32'h83987f11;
    ram_cell[     765] = 32'hc15cdb04;
    ram_cell[     766] = 32'hc8da299b;
    ram_cell[     767] = 32'hfa643b4c;
end

endmodule

